// nios.v

// Generated using ACDS version 13.0 156 at 2018.08.05.10:32:19

`timescale 1 ps / 1 ps
module nios (
		output wire [0:0]  read_n_to_the_ext_flash,                        // flash_ssram_tristate_bridge_bridge_0_out.read_n_to_the_ext_flash
		output wire [0:0]  select_n_to_the_ext_flash,                      //                                         .select_n_to_the_ext_flash
		output wire [25:0] flash_ssram_tristate_bridge_address,            //                                         .flash_ssram_tristate_bridge_address
		output wire [0:0]  bwe_n_to_the_ssram,                             //                                         .bwe_n_to_the_ssram
		output wire [0:0]  reset_n_to_the_ssram,                           //                                         .reset_n_to_the_ssram
		output wire [0:0]  chipenable1_n_to_the_ssram,                     //                                         .chipenable1_n_to_the_ssram
		output wire [3:0]  bw_n_to_the_ssram,                              //                                         .bw_n_to_the_ssram
		output wire [0:0]  outputenable_n_to_the_ssram,                    //                                         .outputenable_n_to_the_ssram
		inout  wire [31:0] flash_ssram_tristate_bridge_data,               //                                         .flash_ssram_tristate_bridge_data
		output wire [0:0]  adsc_n_to_the_ssram,                            //                                         .adsc_n_to_the_ssram
		output wire [19:0] address_to_the_ssram,                           //                                         .address_to_the_ssram
		output wire [0:0]  write_n_to_the_ext_flash,                       //                                         .write_n_to_the_ext_flash
		input  wire        clk,                                            //                               clk_clk_in.clk
		input  wire        clk_125,                                        //                           clk_125_clk_in.clk
		output wire        pll_c0_out,                                     //                               c0_out_clk.clk
		output wire        pll_c2_out,                                     //                               c2_out_clk.clk
		input  wire [3:0]  button_pio_external_connection_export,          //           button_pio_external_connection.export
		output wire [7:0]  led_pio_external_connection_export,             //              led_pio_external_connection.export
		output wire        lcd_display_external_RS,                        //                     lcd_display_external.RS
		output wire        lcd_display_external_RW,                        //                                         .RW
		inout  wire [7:0]  lcd_display_external_data,                      //                                         .data
		output wire        lcd_display_external_E,                         //                                         .E
		output wire [15:0] seven_seg_pio_external_connection_export,       //        seven_seg_pio_external_connection.export
		output wire        ddr2_top_external_connection_local_refresh_ack, //             ddr2_top_external_connection.local_refresh_ack
		output wire        ddr2_top_external_connection_local_init_done,   //                                         .local_init_done
		output wire        ddr2_top_external_connection_reset_phy_clk_n,   //                                         .reset_phy_clk_n
		output wire [0:0]  ddr2_top_memory_mem_odt,                        //                          ddr2_top_memory.mem_odt
		inout  wire [0:0]  ddr2_top_memory_mem_clk,                        //                                         .mem_clk
		inout  wire [0:0]  ddr2_top_memory_mem_clk_n,                      //                                         .mem_clk_n
		output wire [0:0]  ddr2_top_memory_mem_cs_n,                       //                                         .mem_cs_n
		output wire [0:0]  ddr2_top_memory_mem_cke,                        //                                         .mem_cke
		output wire [12:0] ddr2_top_memory_mem_addr,                       //                                         .mem_addr
		output wire [1:0]  ddr2_top_memory_mem_ba,                         //                                         .mem_ba
		output wire        ddr2_top_memory_mem_ras_n,                      //                                         .mem_ras_n
		output wire        ddr2_top_memory_mem_cas_n,                      //                                         .mem_cas_n
		output wire        ddr2_top_memory_mem_we_n,                       //                                         .mem_we_n
		inout  wire [31:0] ddr2_top_memory_mem_dq,                         //                                         .mem_dq
		inout  wire [3:0]  ddr2_top_memory_mem_dqs,                        //                                         .mem_dqs
		output wire [3:0]  ddr2_top_memory_mem_dm,                         //                                         .mem_dm
		output wire        ddr2_top_auxfull_clk,                           //                         ddr2_top_auxfull.clk
		output wire        ddr2_top_auxhalf_clk,                           //                         ddr2_top_auxhalf.clk
		output wire        sysclk_top_out_clk_clk,                         //                       sysclk_top_out_clk.clk
		output wire        ddr2_bot_external_connection_local_refresh_ack, //             ddr2_bot_external_connection.local_refresh_ack
		output wire        ddr2_bot_external_connection_local_init_done,   //                                         .local_init_done
		output wire        ddr2_bot_external_connection_reset_phy_clk_n,   //                                         .reset_phy_clk_n
		output wire [0:0]  ddr2_bot_memory_mem_odt,                        //                          ddr2_bot_memory.mem_odt
		inout  wire [0:0]  ddr2_bot_memory_mem_clk,                        //                                         .mem_clk
		inout  wire [0:0]  ddr2_bot_memory_mem_clk_n,                      //                                         .mem_clk_n
		output wire [0:0]  ddr2_bot_memory_mem_cs_n,                       //                                         .mem_cs_n
		output wire [0:0]  ddr2_bot_memory_mem_cke,                        //                                         .mem_cke
		output wire [12:0] ddr2_bot_memory_mem_addr,                       //                                         .mem_addr
		output wire [1:0]  ddr2_bot_memory_mem_ba,                         //                                         .mem_ba
		output wire        ddr2_bot_memory_mem_ras_n,                      //                                         .mem_ras_n
		output wire        ddr2_bot_memory_mem_cas_n,                      //                                         .mem_cas_n
		output wire        ddr2_bot_memory_mem_we_n,                       //                                         .mem_we_n
		inout  wire [31:0] ddr2_bot_memory_mem_dq,                         //                                         .mem_dq
		inout  wire [3:0]  ddr2_bot_memory_mem_dqs,                        //                                         .mem_dqs
		output wire [3:0]  ddr2_bot_memory_mem_dm,                         //                                         .mem_dm
		output wire        sysclk_bot_out_clk_clk,                         //                       sysclk_bot_out_clk.clk
		input  wire        merged_resets_in_reset_reset_n                  //                   merged_resets_in_reset.reset_n
	);

	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out;                              // flash_ssram_tristate_bridge_pinSharer_0:select_n_to_the_ext_flash -> flash_ssram_tristate_bridge_bridge_0:tcs_select_n_to_the_ext_flash
	wire          flash_ssram_tristate_bridge_pinsharer_0_tcm_grant;                                                      // flash_ssram_tristate_bridge_bridge_0:grant -> flash_ssram_tristate_bridge_pinSharer_0:grant
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_outputenable_n_to_the_ssram_out;                            // flash_ssram_tristate_bridge_pinSharer_0:outputenable_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_outputenable_n_to_the_ssram
	wire   [31:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_in;                        // flash_ssram_tristate_bridge_bridge_0:tcs_flash_ssram_tristate_bridge_data_in -> flash_ssram_tristate_bridge_pinSharer_0:flash_ssram_tristate_bridge_data_in
	wire   [25:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_address_out;                    // flash_ssram_tristate_bridge_pinSharer_0:flash_ssram_tristate_bridge_address -> flash_ssram_tristate_bridge_bridge_0:tcs_flash_ssram_tristate_bridge_address
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out;                                // flash_ssram_tristate_bridge_pinSharer_0:read_n_to_the_ext_flash -> flash_ssram_tristate_bridge_bridge_0:tcs_read_n_to_the_ext_flash
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_adsc_n_to_the_ssram_out;                                    // flash_ssram_tristate_bridge_pinSharer_0:adsc_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_adsc_n_to_the_ssram
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out;                               // flash_ssram_tristate_bridge_pinSharer_0:write_n_to_the_ext_flash -> flash_ssram_tristate_bridge_bridge_0:tcs_write_n_to_the_ext_flash
	wire   [19:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_address_to_the_ssram_out;                                   // flash_ssram_tristate_bridge_pinSharer_0:address_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_address_to_the_ssram
	wire          flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_outen;                     // flash_ssram_tristate_bridge_pinSharer_0:flash_ssram_tristate_bridge_data_outen -> flash_ssram_tristate_bridge_bridge_0:tcs_flash_ssram_tristate_bridge_data_outen
	wire   [31:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_out;                       // flash_ssram_tristate_bridge_pinSharer_0:flash_ssram_tristate_bridge_data -> flash_ssram_tristate_bridge_bridge_0:tcs_flash_ssram_tristate_bridge_data
	wire          flash_ssram_tristate_bridge_pinsharer_0_tcm_request;                                                    // flash_ssram_tristate_bridge_pinSharer_0:request -> flash_ssram_tristate_bridge_bridge_0:request
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_bwe_n_to_the_ssram_out;                                     // flash_ssram_tristate_bridge_pinSharer_0:bwe_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_bwe_n_to_the_ssram
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_reset_n_to_the_ssram_out;                                   // flash_ssram_tristate_bridge_pinSharer_0:reset_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_reset_n_to_the_ssram
	wire    [0:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_chipenable1_n_to_the_ssram_out;                             // flash_ssram_tristate_bridge_pinSharer_0:chipenable1_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_chipenable1_n_to_the_ssram
	wire    [3:0] flash_ssram_tristate_bridge_pinsharer_0_tcm_bw_n_to_the_ssram_out;                                      // flash_ssram_tristate_bridge_pinSharer_0:bw_n_to_the_ssram -> flash_ssram_tristate_bridge_bridge_0:tcs_bw_n_to_the_ssram
	wire          ssram_tcm_chipselect_n_out;                                                                             // ssram:tcm_chipselect_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_chipselect_n_out
	wire          ssram_tcm_grant;                                                                                        // flash_ssram_tristate_bridge_pinSharer_0:tcs0_grant -> ssram:tcm_grant
	wire          ssram_tcm_data_outen;                                                                                   // ssram:tcm_data_outen -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_data_outen
	wire          ssram_tcm_reset_n_out;                                                                                  // ssram:tcm_reset_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_reset_n_out
	wire          ssram_tcm_outputenable_n_out;                                                                           // ssram:tcm_outputenable_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_outputenable_n_out
	wire          ssram_tcm_request;                                                                                      // ssram:tcm_request -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_request
	wire   [31:0] ssram_tcm_data_out;                                                                                     // ssram:tcm_data_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_data_out
	wire          ssram_tcm_write_n_out;                                                                                  // ssram:tcm_write_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_write_n_out
	wire   [19:0] ssram_tcm_address_out;                                                                                  // ssram:tcm_address_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_address_out
	wire   [31:0] ssram_tcm_data_in;                                                                                      // flash_ssram_tristate_bridge_pinSharer_0:tcs0_data_in -> ssram:tcm_data_in
	wire          ssram_tcm_begintransfer_n_out;                                                                          // ssram:tcm_begintransfer_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_begintransfer_n_out
	wire    [3:0] ssram_tcm_byteenable_n_out;                                                                             // ssram:tcm_byteenable_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs0_byteenable_n_out
	wire          ext_flash_tcm_chipselect_n_out;                                                                         // ext_flash:tcm_chipselect_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_chipselect_n_out
	wire          ext_flash_tcm_grant;                                                                                    // flash_ssram_tristate_bridge_pinSharer_0:tcs1_grant -> ext_flash:tcm_grant
	wire          ext_flash_tcm_data_outen;                                                                               // ext_flash:tcm_data_outen -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_data_outen
	wire          ext_flash_tcm_request;                                                                                  // ext_flash:tcm_request -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_request
	wire   [15:0] ext_flash_tcm_data_out;                                                                                 // ext_flash:tcm_data_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_data_out
	wire          ext_flash_tcm_write_n_out;                                                                              // ext_flash:tcm_write_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_write_n_out
	wire   [25:0] ext_flash_tcm_address_out;                                                                              // ext_flash:tcm_address_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_address_out
	wire   [15:0] ext_flash_tcm_data_in;                                                                                  // flash_ssram_tristate_bridge_pinSharer_0:tcs1_data_in -> ext_flash:tcm_data_in
	wire          ext_flash_tcm_read_n_out;                                                                               // ext_flash:tcm_read_n_out -> flash_ssram_tristate_bridge_pinSharer_0:tcs1_read_n_out
	wire    [2:0] fir_dma_write_master_burstcount;                                                                        // fir_dma:write_master_burstcount -> fir_dma_write_master_translator:av_burstcount
	wire          fir_dma_write_master_waitrequest;                                                                       // fir_dma_write_master_translator:av_waitrequest -> fir_dma:write_master_waitrequest
	wire   [31:0] fir_dma_write_master_writedata;                                                                         // fir_dma:write_master_writedata -> fir_dma_write_master_translator:av_writedata
	wire   [31:0] fir_dma_write_master_address;                                                                           // fir_dma:write_master_address -> fir_dma_write_master_translator:av_address
	wire          fir_dma_write_master_write;                                                                             // fir_dma:write_master_write -> fir_dma_write_master_translator:av_write
	wire    [3:0] fir_dma_write_master_byteenable;                                                                        // fir_dma:write_master_byteenable -> fir_dma_write_master_translator:av_byteenable
	wire    [0:0] ddr2_top_clock_bridge_m0_burstcount;                                                                    // ddr2_top_clock_bridge:m0_burstcount -> ddr2_top_clock_bridge_m0_translator:av_burstcount
	wire          ddr2_top_clock_bridge_m0_waitrequest;                                                                   // ddr2_top_clock_bridge_m0_translator:av_waitrequest -> ddr2_top_clock_bridge:m0_waitrequest
	wire   [26:0] ddr2_top_clock_bridge_m0_address;                                                                       // ddr2_top_clock_bridge:m0_address -> ddr2_top_clock_bridge_m0_translator:av_address
	wire  [127:0] ddr2_top_clock_bridge_m0_writedata;                                                                     // ddr2_top_clock_bridge:m0_writedata -> ddr2_top_clock_bridge_m0_translator:av_writedata
	wire          ddr2_top_clock_bridge_m0_write;                                                                         // ddr2_top_clock_bridge:m0_write -> ddr2_top_clock_bridge_m0_translator:av_write
	wire          ddr2_top_clock_bridge_m0_read;                                                                          // ddr2_top_clock_bridge:m0_read -> ddr2_top_clock_bridge_m0_translator:av_read
	wire  [127:0] ddr2_top_clock_bridge_m0_readdata;                                                                      // ddr2_top_clock_bridge_m0_translator:av_readdata -> ddr2_top_clock_bridge:m0_readdata
	wire          ddr2_top_clock_bridge_m0_debugaccess;                                                                   // ddr2_top_clock_bridge:m0_debugaccess -> ddr2_top_clock_bridge_m0_translator:av_debugaccess
	wire   [15:0] ddr2_top_clock_bridge_m0_byteenable;                                                                    // ddr2_top_clock_bridge:m0_byteenable -> ddr2_top_clock_bridge_m0_translator:av_byteenable
	wire          ddr2_top_clock_bridge_m0_readdatavalid;                                                                 // ddr2_top_clock_bridge_m0_translator:av_readdatavalid -> ddr2_top_clock_bridge:m0_readdatavalid
	wire          ddr2_top_s1_translator_avalon_anti_slave_0_waitrequest;                                                 // ddr2_top:local_ready -> ddr2_top_s1_translator:av_waitrequest
	wire    [2:0] ddr2_top_s1_translator_avalon_anti_slave_0_burstcount;                                                  // ddr2_top_s1_translator:av_burstcount -> ddr2_top:local_size
	wire   [63:0] ddr2_top_s1_translator_avalon_anti_slave_0_writedata;                                                   // ddr2_top_s1_translator:av_writedata -> ddr2_top:local_wdata
	wire   [23:0] ddr2_top_s1_translator_avalon_anti_slave_0_address;                                                     // ddr2_top_s1_translator:av_address -> ddr2_top:local_address
	wire          ddr2_top_s1_translator_avalon_anti_slave_0_write;                                                       // ddr2_top_s1_translator:av_write -> ddr2_top:local_write_req
	wire          ddr2_top_s1_translator_avalon_anti_slave_0_beginbursttransfer;                                          // ddr2_top_s1_translator:av_beginbursttransfer -> ddr2_top:local_burstbegin
	wire          ddr2_top_s1_translator_avalon_anti_slave_0_read;                                                        // ddr2_top_s1_translator:av_read -> ddr2_top:local_read_req
	wire   [63:0] ddr2_top_s1_translator_avalon_anti_slave_0_readdata;                                                    // ddr2_top:local_rdata -> ddr2_top_s1_translator:av_readdata
	wire          ddr2_top_s1_translator_avalon_anti_slave_0_readdatavalid;                                               // ddr2_top:local_rdata_valid -> ddr2_top_s1_translator:av_readdatavalid
	wire    [7:0] ddr2_top_s1_translator_avalon_anti_slave_0_byteenable;                                                  // ddr2_top_s1_translator:av_byteenable -> ddr2_top:local_be
	wire          ddr2_top_reset_request_n_reset;                                                                         // ddr2_top:reset_request_n -> [cmd_xbar_mux:reset, crosser:out_reset, crosser_001:in_reset, ddr2_top_s1_translator:reset, ddr2_top_s1_translator_avalon_universal_slave_0_agent:reset, ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, rsp_xbar_demux:reset, rst_controller:reset_in2, rst_controller_002:reset_in2, rst_controller_003:reset_in2, rst_controller_004:reset_in2, rst_controller_005:reset_in2, rst_controller_006:reset_in1]
	wire          fir_dma_read_master_waitrequest;                                                                        // fir_dma_read_master_translator:av_waitrequest -> fir_dma:read_master_waitrequest
	wire   [31:0] fir_dma_read_master_address;                                                                            // fir_dma:read_master_address -> fir_dma_read_master_translator:av_address
	wire          fir_dma_read_master_read;                                                                               // fir_dma:read_master_read -> fir_dma_read_master_translator:av_read
	wire   [31:0] fir_dma_read_master_readdata;                                                                           // fir_dma_read_master_translator:av_readdata -> fir_dma:read_master_readdata
	wire          fir_dma_read_master_readdatavalid;                                                                      // fir_dma_read_master_translator:av_readdatavalid -> fir_dma:read_master_readdatavalid
	wire    [3:0] fir_dma_read_master_byteenable;                                                                         // fir_dma:read_master_byteenable -> fir_dma_read_master_translator:av_byteenable
	wire          cpu_data_master_waitrequest;                                                                            // cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                                                              // cpu:d_writedata -> cpu_data_master_translator:av_writedata
	wire   [29:0] cpu_data_master_address;                                                                                // cpu:d_address -> cpu_data_master_translator:av_address
	wire          cpu_data_master_write;                                                                                  // cpu:d_write -> cpu_data_master_translator:av_write
	wire          cpu_data_master_read;                                                                                   // cpu:d_read -> cpu_data_master_translator:av_read
	wire   [31:0] cpu_data_master_readdata;                                                                               // cpu_data_master_translator:av_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                                                            // cpu:jtag_debug_module_debugaccess_to_roms -> cpu_data_master_translator:av_debugaccess
	wire          cpu_data_master_readdatavalid;                                                                          // cpu_data_master_translator:av_readdatavalid -> cpu:d_readdatavalid
	wire    [3:0] cpu_data_master_byteenable;                                                                             // cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	wire          cpu_instruction_master_waitrequest;                                                                     // cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	wire   [29:0] cpu_instruction_master_address;                                                                         // cpu:i_address -> cpu_instruction_master_translator:av_address
	wire          cpu_instruction_master_read;                                                                            // cpu:i_read -> cpu_instruction_master_translator:av_read
	wire   [31:0] cpu_instruction_master_readdata;                                                                        // cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                                                                   // cpu_instruction_master_translator:av_readdatavalid -> cpu:i_readdatavalid
	wire          dma_0_read_master_waitrequest;                                                                          // dma_0_read_master_translator:av_waitrequest -> dma_0:read_waitrequest
	wire   [29:0] dma_0_read_master_address;                                                                              // dma_0:read_address -> dma_0_read_master_translator:av_address
	wire          dma_0_read_master_chipselect;                                                                           // dma_0:read_chipselect -> dma_0_read_master_translator:av_chipselect
	wire          dma_0_read_master_read;                                                                                 // dma_0:read_read_n -> dma_0_read_master_translator:av_read
	wire  [127:0] dma_0_read_master_readdata;                                                                             // dma_0_read_master_translator:av_readdata -> dma_0:read_readdata
	wire          dma_0_read_master_readdatavalid;                                                                        // dma_0_read_master_translator:av_readdatavalid -> dma_0:read_readdatavalid
	wire          dma_0_write_master_waitrequest;                                                                         // dma_0_write_master_translator:av_waitrequest -> dma_0:write_waitrequest
	wire  [127:0] dma_0_write_master_writedata;                                                                           // dma_0:write_writedata -> dma_0_write_master_translator:av_writedata
	wire   [28:0] dma_0_write_master_address;                                                                             // dma_0:write_address -> dma_0_write_master_translator:av_address
	wire          dma_0_write_master_chipselect;                                                                          // dma_0:write_chipselect -> dma_0_write_master_translator:av_chipselect
	wire          dma_0_write_master_write;                                                                               // dma_0:write_write_n -> dma_0_write_master_translator:av_write
	wire   [15:0] dma_0_write_master_byteenable;                                                                          // dma_0:write_byteenable -> dma_0_write_master_translator:av_byteenable
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                              // flash_ssram_pipeline_bridge:s0_waitrequest -> flash_ssram_pipeline_bridge_s0_translator:av_waitrequest
	wire    [0:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_burstcount;                               // flash_ssram_pipeline_bridge_s0_translator:av_burstcount -> flash_ssram_pipeline_bridge:s0_burstcount
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_writedata;                                // flash_ssram_pipeline_bridge_s0_translator:av_writedata -> flash_ssram_pipeline_bridge:s0_writedata
	wire   [26:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_address;                                  // flash_ssram_pipeline_bridge_s0_translator:av_address -> flash_ssram_pipeline_bridge:s0_address
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_write;                                    // flash_ssram_pipeline_bridge_s0_translator:av_write -> flash_ssram_pipeline_bridge:s0_write
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_read;                                     // flash_ssram_pipeline_bridge_s0_translator:av_read -> flash_ssram_pipeline_bridge:s0_read
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdata;                                 // flash_ssram_pipeline_bridge:s0_readdata -> flash_ssram_pipeline_bridge_s0_translator:av_readdata
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                              // flash_ssram_pipeline_bridge_s0_translator:av_debugaccess -> flash_ssram_pipeline_bridge:s0_debugaccess
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                            // flash_ssram_pipeline_bridge:s0_readdatavalid -> flash_ssram_pipeline_bridge_s0_translator:av_readdatavalid
	wire    [3:0] flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_byteenable;                               // flash_ssram_pipeline_bridge_s0_translator:av_byteenable -> flash_ssram_pipeline_bridge:s0_byteenable
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                   // slow_peripheral_bridge:s0_waitrequest -> slow_peripheral_bridge_s0_translator:av_waitrequest
	wire    [0:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                    // slow_peripheral_bridge_s0_translator:av_burstcount -> slow_peripheral_bridge:s0_burstcount
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata;                                     // slow_peripheral_bridge_s0_translator:av_writedata -> slow_peripheral_bridge:s0_writedata
	wire    [9:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address;                                       // slow_peripheral_bridge_s0_translator:av_address -> slow_peripheral_bridge:s0_address
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write;                                         // slow_peripheral_bridge_s0_translator:av_write -> slow_peripheral_bridge:s0_write
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read;                                          // slow_peripheral_bridge_s0_translator:av_read -> slow_peripheral_bridge:s0_read
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata;                                      // slow_peripheral_bridge:s0_readdata -> slow_peripheral_bridge_s0_translator:av_readdata
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                   // slow_peripheral_bridge_s0_translator:av_debugaccess -> slow_peripheral_bridge:s0_debugaccess
	wire          slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                 // slow_peripheral_bridge:s0_readdatavalid -> slow_peripheral_bridge_s0_translator:av_readdatavalid
	wire    [3:0] slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                    // slow_peripheral_bridge_s0_translator:av_byteenable -> slow_peripheral_bridge:s0_byteenable
	wire          ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                    // ddr2_top_clock_bridge:s0_waitrequest -> ddr2_top_clock_bridge_s0_translator:av_waitrequest
	wire    [0:0] ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                     // ddr2_top_clock_bridge_s0_translator:av_burstcount -> ddr2_top_clock_bridge:s0_burstcount
	wire  [127:0] ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_writedata;                                      // ddr2_top_clock_bridge_s0_translator:av_writedata -> ddr2_top_clock_bridge:s0_writedata
	wire   [26:0] ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_address;                                        // ddr2_top_clock_bridge_s0_translator:av_address -> ddr2_top_clock_bridge:s0_address
	wire          ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_write;                                          // ddr2_top_clock_bridge_s0_translator:av_write -> ddr2_top_clock_bridge:s0_write
	wire          ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_read;                                           // ddr2_top_clock_bridge_s0_translator:av_read -> ddr2_top_clock_bridge:s0_read
	wire  [127:0] ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_readdata;                                       // ddr2_top_clock_bridge:s0_readdata -> ddr2_top_clock_bridge_s0_translator:av_readdata
	wire          ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                    // ddr2_top_clock_bridge_s0_translator:av_debugaccess -> ddr2_top_clock_bridge:s0_debugaccess
	wire          ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                  // ddr2_top_clock_bridge:s0_readdatavalid -> ddr2_top_clock_bridge_s0_translator:av_readdatavalid
	wire   [15:0] ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                     // ddr2_top_clock_bridge_s0_translator:av_byteenable -> ddr2_top_clock_bridge:s0_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest;                                       // cpu:jtag_debug_module_waitrequest -> cpu_jtag_debug_module_translator:av_waitrequest
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                                         // cpu_jtag_debug_module_translator:av_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_address;                                           // cpu_jtag_debug_module_translator:av_address -> cpu:jtag_debug_module_address
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_write;                                             // cpu_jtag_debug_module_translator:av_write -> cpu:jtag_debug_module_write
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_read;                                              // cpu_jtag_debug_module_translator:av_read -> cpu:jtag_debug_module_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                                          // cpu:jtag_debug_module_readdata -> cpu_jtag_debug_module_translator:av_readdata
	wire          cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                                       // cpu_jtag_debug_module_translator:av_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                                        // cpu_jtag_debug_module_translator:av_byteenable -> cpu:jtag_debug_module_byteenable
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest;                                    // ddr2_bot_clock_bridge:s0_waitrequest -> ddr2_bot_clock_bridge_s0_translator:av_waitrequest
	wire    [0:0] ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount;                                     // ddr2_bot_clock_bridge_s0_translator:av_burstcount -> ddr2_bot_clock_bridge:s0_burstcount
	wire  [127:0] ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_writedata;                                      // ddr2_bot_clock_bridge_s0_translator:av_writedata -> ddr2_bot_clock_bridge:s0_writedata
	wire   [26:0] ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_address;                                        // ddr2_bot_clock_bridge_s0_translator:av_address -> ddr2_bot_clock_bridge:s0_address
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_write;                                          // ddr2_bot_clock_bridge_s0_translator:av_write -> ddr2_bot_clock_bridge:s0_write
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_read;                                           // ddr2_bot_clock_bridge_s0_translator:av_read -> ddr2_bot_clock_bridge:s0_read
	wire  [127:0] ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_readdata;                                       // ddr2_bot_clock_bridge:s0_readdata -> ddr2_bot_clock_bridge_s0_translator:av_readdata
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess;                                    // ddr2_bot_clock_bridge_s0_translator:av_debugaccess -> ddr2_bot_clock_bridge:s0_debugaccess
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid;                                  // ddr2_bot_clock_bridge:s0_readdatavalid -> ddr2_bot_clock_bridge_s0_translator:av_readdatavalid
	wire   [15:0] ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable;                                     // ddr2_bot_clock_bridge_s0_translator:av_byteenable -> ddr2_bot_clock_bridge:s0_byteenable
	wire   [31:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata;                                      // dma_0_control_port_slave_translator:av_writedata -> dma_0:dma_ctl_writedata
	wire    [2:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_address;                                        // dma_0_control_port_slave_translator:av_address -> dma_0:dma_ctl_address
	wire          dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect;                                     // dma_0_control_port_slave_translator:av_chipselect -> dma_0:dma_ctl_chipselect
	wire          dma_0_control_port_slave_translator_avalon_anti_slave_0_write;                                          // dma_0_control_port_slave_translator:av_write -> dma_0:dma_ctl_write_n
	wire   [31:0] dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata;                                       // dma_0:dma_ctl_readdata -> dma_0_control_port_slave_translator:av_readdata
	wire    [0:0] slow_peripheral_bridge_m0_burstcount;                                                                   // slow_peripheral_bridge:m0_burstcount -> slow_peripheral_bridge_m0_translator:av_burstcount
	wire          slow_peripheral_bridge_m0_waitrequest;                                                                  // slow_peripheral_bridge_m0_translator:av_waitrequest -> slow_peripheral_bridge:m0_waitrequest
	wire    [9:0] slow_peripheral_bridge_m0_address;                                                                      // slow_peripheral_bridge:m0_address -> slow_peripheral_bridge_m0_translator:av_address
	wire   [31:0] slow_peripheral_bridge_m0_writedata;                                                                    // slow_peripheral_bridge:m0_writedata -> slow_peripheral_bridge_m0_translator:av_writedata
	wire          slow_peripheral_bridge_m0_write;                                                                        // slow_peripheral_bridge:m0_write -> slow_peripheral_bridge_m0_translator:av_write
	wire          slow_peripheral_bridge_m0_read;                                                                         // slow_peripheral_bridge:m0_read -> slow_peripheral_bridge_m0_translator:av_read
	wire   [31:0] slow_peripheral_bridge_m0_readdata;                                                                     // slow_peripheral_bridge_m0_translator:av_readdata -> slow_peripheral_bridge:m0_readdata
	wire          slow_peripheral_bridge_m0_debugaccess;                                                                  // slow_peripheral_bridge:m0_debugaccess -> slow_peripheral_bridge_m0_translator:av_debugaccess
	wire    [3:0] slow_peripheral_bridge_m0_byteenable;                                                                   // slow_peripheral_bridge:m0_byteenable -> slow_peripheral_bridge_m0_translator:av_byteenable
	wire          slow_peripheral_bridge_m0_readdatavalid;                                                                // slow_peripheral_bridge_m0_translator:av_readdatavalid -> slow_peripheral_bridge:m0_readdatavalid
	wire   [15:0] high_res_timer_s1_translator_avalon_anti_slave_0_writedata;                                             // high_res_timer_s1_translator:av_writedata -> high_res_timer:writedata
	wire    [2:0] high_res_timer_s1_translator_avalon_anti_slave_0_address;                                               // high_res_timer_s1_translator:av_address -> high_res_timer:address
	wire          high_res_timer_s1_translator_avalon_anti_slave_0_chipselect;                                            // high_res_timer_s1_translator:av_chipselect -> high_res_timer:chipselect
	wire          high_res_timer_s1_translator_avalon_anti_slave_0_write;                                                 // high_res_timer_s1_translator:av_write -> high_res_timer:write_n
	wire   [15:0] high_res_timer_s1_translator_avalon_anti_slave_0_readdata;                                              // high_res_timer:readdata -> high_res_timer_s1_translator:av_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                                 // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                   // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                     // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                                  // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                       // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                        // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                    // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire   [31:0] performance_counter_control_slave_translator_avalon_anti_slave_0_writedata;                             // performance_counter_control_slave_translator:av_writedata -> performance_counter:writedata
	wire    [2:0] performance_counter_control_slave_translator_avalon_anti_slave_0_address;                               // performance_counter_control_slave_translator:av_address -> performance_counter:address
	wire          performance_counter_control_slave_translator_avalon_anti_slave_0_write;                                 // performance_counter_control_slave_translator:av_write -> performance_counter:write
	wire   [31:0] performance_counter_control_slave_translator_avalon_anti_slave_0_readdata;                              // performance_counter:readdata -> performance_counter_control_slave_translator:av_readdata
	wire          performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer;                         // performance_counter_control_slave_translator:av_begintransfer -> performance_counter:begintransfer
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata;                                              // sys_clk_timer_s1_translator:av_writedata -> sys_clk_timer:writedata
	wire    [2:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_address;                                                // sys_clk_timer_s1_translator:av_address -> sys_clk_timer:address
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect;                                             // sys_clk_timer_s1_translator:av_chipselect -> sys_clk_timer:chipselect
	wire          sys_clk_timer_s1_translator_avalon_anti_slave_0_write;                                                  // sys_clk_timer_s1_translator:av_write -> sys_clk_timer:write_n
	wire   [15:0] sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata;                                               // sys_clk_timer:readdata -> sys_clk_timer_s1_translator:av_readdata
	wire    [0:0] sysid_control_slave_translator_avalon_anti_slave_0_address;                                             // sysid_control_slave_translator:av_address -> sysid:address
	wire   [31:0] sysid_control_slave_translator_avalon_anti_slave_0_readdata;                                            // sysid:readdata -> sysid_control_slave_translator:av_readdata
	wire   [31:0] fir_dma_control_translator_avalon_anti_slave_0_writedata;                                               // fir_dma_control_translator:av_writedata -> fir_dma:slave_writedata
	wire    [2:0] fir_dma_control_translator_avalon_anti_slave_0_address;                                                 // fir_dma_control_translator:av_address -> fir_dma:slave_address
	wire          fir_dma_control_translator_avalon_anti_slave_0_write;                                                   // fir_dma_control_translator:av_write -> fir_dma:slave_write
	wire          fir_dma_control_translator_avalon_anti_slave_0_read;                                                    // fir_dma_control_translator:av_read -> fir_dma:slave_read
	wire   [31:0] fir_dma_control_translator_avalon_anti_slave_0_readdata;                                                // fir_dma:slave_readdata -> fir_dma_control_translator:av_readdata
	wire    [3:0] fir_dma_control_translator_avalon_anti_slave_0_byteenable;                                              // fir_dma_control_translator:av_byteenable -> fir_dma:slave_byteenable
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_writedata;                                                 // pll_pll_slave_translator:av_writedata -> pll:writedata
	wire    [1:0] pll_pll_slave_translator_avalon_anti_slave_0_address;                                                   // pll_pll_slave_translator:av_address -> pll:address
	wire          pll_pll_slave_translator_avalon_anti_slave_0_write;                                                     // pll_pll_slave_translator:av_write -> pll:write
	wire          pll_pll_slave_translator_avalon_anti_slave_0_read;                                                      // pll_pll_slave_translator:av_read -> pll:read
	wire   [31:0] pll_pll_slave_translator_avalon_anti_slave_0_readdata;                                                  // pll:readdata -> pll_pll_slave_translator:av_readdata
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_writedata;                                                 // button_pio_s1_translator:av_writedata -> button_pio:writedata
	wire    [1:0] button_pio_s1_translator_avalon_anti_slave_0_address;                                                   // button_pio_s1_translator:av_address -> button_pio:address
	wire          button_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                // button_pio_s1_translator:av_chipselect -> button_pio:chipselect
	wire          button_pio_s1_translator_avalon_anti_slave_0_write;                                                     // button_pio_s1_translator:av_write -> button_pio:write_n
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_readdata;                                                  // button_pio:readdata -> button_pio_s1_translator:av_readdata
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_writedata;                                                    // led_pio_s1_translator:av_writedata -> led_pio:writedata
	wire    [1:0] led_pio_s1_translator_avalon_anti_slave_0_address;                                                      // led_pio_s1_translator:av_address -> led_pio:address
	wire          led_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                   // led_pio_s1_translator:av_chipselect -> led_pio:chipselect
	wire          led_pio_s1_translator_avalon_anti_slave_0_write;                                                        // led_pio_s1_translator:av_write -> led_pio:write_n
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_readdata;                                                     // led_pio:readdata -> led_pio_s1_translator:av_readdata
	wire    [7:0] lcd_display_control_slave_translator_avalon_anti_slave_0_writedata;                                     // lcd_display_control_slave_translator:av_writedata -> lcd_display:writedata
	wire    [1:0] lcd_display_control_slave_translator_avalon_anti_slave_0_address;                                       // lcd_display_control_slave_translator:av_address -> lcd_display:address
	wire          lcd_display_control_slave_translator_avalon_anti_slave_0_write;                                         // lcd_display_control_slave_translator:av_write -> lcd_display:write
	wire          lcd_display_control_slave_translator_avalon_anti_slave_0_read;                                          // lcd_display_control_slave_translator:av_read -> lcd_display:read
	wire    [7:0] lcd_display_control_slave_translator_avalon_anti_slave_0_readdata;                                      // lcd_display:readdata -> lcd_display_control_slave_translator:av_readdata
	wire          lcd_display_control_slave_translator_avalon_anti_slave_0_begintransfer;                                 // lcd_display_control_slave_translator:av_begintransfer -> lcd_display:begintransfer
	wire   [31:0] seven_seg_pio_s1_translator_avalon_anti_slave_0_writedata;                                              // seven_seg_pio_s1_translator:av_writedata -> seven_seg_pio:writedata
	wire    [1:0] seven_seg_pio_s1_translator_avalon_anti_slave_0_address;                                                // seven_seg_pio_s1_translator:av_address -> seven_seg_pio:address
	wire          seven_seg_pio_s1_translator_avalon_anti_slave_0_chipselect;                                             // seven_seg_pio_s1_translator:av_chipselect -> seven_seg_pio:chipselect
	wire          seven_seg_pio_s1_translator_avalon_anti_slave_0_write;                                                  // seven_seg_pio_s1_translator:av_write -> seven_seg_pio:write_n
	wire   [31:0] seven_seg_pio_s1_translator_avalon_anti_slave_0_readdata;                                               // seven_seg_pio:readdata -> seven_seg_pio_s1_translator:av_readdata
	wire    [0:0] flash_ssram_pipeline_bridge_m0_burstcount;                                                              // flash_ssram_pipeline_bridge:m0_burstcount -> flash_ssram_pipeline_bridge_m0_translator:av_burstcount
	wire          flash_ssram_pipeline_bridge_m0_waitrequest;                                                             // flash_ssram_pipeline_bridge_m0_translator:av_waitrequest -> flash_ssram_pipeline_bridge:m0_waitrequest
	wire   [26:0] flash_ssram_pipeline_bridge_m0_address;                                                                 // flash_ssram_pipeline_bridge:m0_address -> flash_ssram_pipeline_bridge_m0_translator:av_address
	wire   [31:0] flash_ssram_pipeline_bridge_m0_writedata;                                                               // flash_ssram_pipeline_bridge:m0_writedata -> flash_ssram_pipeline_bridge_m0_translator:av_writedata
	wire          flash_ssram_pipeline_bridge_m0_write;                                                                   // flash_ssram_pipeline_bridge:m0_write -> flash_ssram_pipeline_bridge_m0_translator:av_write
	wire          flash_ssram_pipeline_bridge_m0_read;                                                                    // flash_ssram_pipeline_bridge:m0_read -> flash_ssram_pipeline_bridge_m0_translator:av_read
	wire   [31:0] flash_ssram_pipeline_bridge_m0_readdata;                                                                // flash_ssram_pipeline_bridge_m0_translator:av_readdata -> flash_ssram_pipeline_bridge:m0_readdata
	wire          flash_ssram_pipeline_bridge_m0_debugaccess;                                                             // flash_ssram_pipeline_bridge:m0_debugaccess -> flash_ssram_pipeline_bridge_m0_translator:av_debugaccess
	wire    [3:0] flash_ssram_pipeline_bridge_m0_byteenable;                                                              // flash_ssram_pipeline_bridge:m0_byteenable -> flash_ssram_pipeline_bridge_m0_translator:av_byteenable
	wire          flash_ssram_pipeline_bridge_m0_readdatavalid;                                                           // flash_ssram_pipeline_bridge_m0_translator:av_readdatavalid -> flash_ssram_pipeline_bridge:m0_readdatavalid
	wire          ssram_uas_translator_avalon_anti_slave_0_waitrequest;                                                   // ssram:uas_waitrequest -> ssram_uas_translator:av_waitrequest
	wire    [2:0] ssram_uas_translator_avalon_anti_slave_0_burstcount;                                                    // ssram_uas_translator:av_burstcount -> ssram:uas_burstcount
	wire   [31:0] ssram_uas_translator_avalon_anti_slave_0_writedata;                                                     // ssram_uas_translator:av_writedata -> ssram:uas_writedata
	wire   [19:0] ssram_uas_translator_avalon_anti_slave_0_address;                                                       // ssram_uas_translator:av_address -> ssram:uas_address
	wire          ssram_uas_translator_avalon_anti_slave_0_lock;                                                          // ssram_uas_translator:av_lock -> ssram:uas_lock
	wire          ssram_uas_translator_avalon_anti_slave_0_write;                                                         // ssram_uas_translator:av_write -> ssram:uas_write
	wire          ssram_uas_translator_avalon_anti_slave_0_read;                                                          // ssram_uas_translator:av_read -> ssram:uas_read
	wire   [31:0] ssram_uas_translator_avalon_anti_slave_0_readdata;                                                      // ssram:uas_readdata -> ssram_uas_translator:av_readdata
	wire          ssram_uas_translator_avalon_anti_slave_0_debugaccess;                                                   // ssram_uas_translator:av_debugaccess -> ssram:uas_debugaccess
	wire          ssram_uas_translator_avalon_anti_slave_0_readdatavalid;                                                 // ssram:uas_readdatavalid -> ssram_uas_translator:av_readdatavalid
	wire    [3:0] ssram_uas_translator_avalon_anti_slave_0_byteenable;                                                    // ssram_uas_translator:av_byteenable -> ssram:uas_byteenable
	wire          ext_flash_uas_translator_avalon_anti_slave_0_waitrequest;                                               // ext_flash:uas_waitrequest -> ext_flash_uas_translator:av_waitrequest
	wire    [1:0] ext_flash_uas_translator_avalon_anti_slave_0_burstcount;                                                // ext_flash_uas_translator:av_burstcount -> ext_flash:uas_burstcount
	wire   [15:0] ext_flash_uas_translator_avalon_anti_slave_0_writedata;                                                 // ext_flash_uas_translator:av_writedata -> ext_flash:uas_writedata
	wire   [25:0] ext_flash_uas_translator_avalon_anti_slave_0_address;                                                   // ext_flash_uas_translator:av_address -> ext_flash:uas_address
	wire          ext_flash_uas_translator_avalon_anti_slave_0_lock;                                                      // ext_flash_uas_translator:av_lock -> ext_flash:uas_lock
	wire          ext_flash_uas_translator_avalon_anti_slave_0_write;                                                     // ext_flash_uas_translator:av_write -> ext_flash:uas_write
	wire          ext_flash_uas_translator_avalon_anti_slave_0_read;                                                      // ext_flash_uas_translator:av_read -> ext_flash:uas_read
	wire   [15:0] ext_flash_uas_translator_avalon_anti_slave_0_readdata;                                                  // ext_flash:uas_readdata -> ext_flash_uas_translator:av_readdata
	wire          ext_flash_uas_translator_avalon_anti_slave_0_debugaccess;                                               // ext_flash_uas_translator:av_debugaccess -> ext_flash:uas_debugaccess
	wire          ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid;                                             // ext_flash:uas_readdatavalid -> ext_flash_uas_translator:av_readdatavalid
	wire    [1:0] ext_flash_uas_translator_avalon_anti_slave_0_byteenable;                                                // ext_flash_uas_translator:av_byteenable -> ext_flash:uas_byteenable
	wire    [0:0] ddr2_bot_clock_bridge_m0_burstcount;                                                                    // ddr2_bot_clock_bridge:m0_burstcount -> ddr2_bot_clock_bridge_m0_translator:av_burstcount
	wire          ddr2_bot_clock_bridge_m0_waitrequest;                                                                   // ddr2_bot_clock_bridge_m0_translator:av_waitrequest -> ddr2_bot_clock_bridge:m0_waitrequest
	wire   [26:0] ddr2_bot_clock_bridge_m0_address;                                                                       // ddr2_bot_clock_bridge:m0_address -> ddr2_bot_clock_bridge_m0_translator:av_address
	wire  [127:0] ddr2_bot_clock_bridge_m0_writedata;                                                                     // ddr2_bot_clock_bridge:m0_writedata -> ddr2_bot_clock_bridge_m0_translator:av_writedata
	wire          ddr2_bot_clock_bridge_m0_write;                                                                         // ddr2_bot_clock_bridge:m0_write -> ddr2_bot_clock_bridge_m0_translator:av_write
	wire          ddr2_bot_clock_bridge_m0_read;                                                                          // ddr2_bot_clock_bridge:m0_read -> ddr2_bot_clock_bridge_m0_translator:av_read
	wire  [127:0] ddr2_bot_clock_bridge_m0_readdata;                                                                      // ddr2_bot_clock_bridge_m0_translator:av_readdata -> ddr2_bot_clock_bridge:m0_readdata
	wire          ddr2_bot_clock_bridge_m0_debugaccess;                                                                   // ddr2_bot_clock_bridge:m0_debugaccess -> ddr2_bot_clock_bridge_m0_translator:av_debugaccess
	wire   [15:0] ddr2_bot_clock_bridge_m0_byteenable;                                                                    // ddr2_bot_clock_bridge:m0_byteenable -> ddr2_bot_clock_bridge_m0_translator:av_byteenable
	wire          ddr2_bot_clock_bridge_m0_readdatavalid;                                                                 // ddr2_bot_clock_bridge_m0_translator:av_readdatavalid -> ddr2_bot_clock_bridge:m0_readdatavalid
	wire          ddr2_bot_s1_translator_avalon_anti_slave_0_waitrequest;                                                 // ddr2_bot:local_ready -> ddr2_bot_s1_translator:av_waitrequest
	wire    [2:0] ddr2_bot_s1_translator_avalon_anti_slave_0_burstcount;                                                  // ddr2_bot_s1_translator:av_burstcount -> ddr2_bot:local_size
	wire   [63:0] ddr2_bot_s1_translator_avalon_anti_slave_0_writedata;                                                   // ddr2_bot_s1_translator:av_writedata -> ddr2_bot:local_wdata
	wire   [23:0] ddr2_bot_s1_translator_avalon_anti_slave_0_address;                                                     // ddr2_bot_s1_translator:av_address -> ddr2_bot:local_address
	wire          ddr2_bot_s1_translator_avalon_anti_slave_0_write;                                                       // ddr2_bot_s1_translator:av_write -> ddr2_bot:local_write_req
	wire          ddr2_bot_s1_translator_avalon_anti_slave_0_beginbursttransfer;                                          // ddr2_bot_s1_translator:av_beginbursttransfer -> ddr2_bot:local_burstbegin
	wire          ddr2_bot_s1_translator_avalon_anti_slave_0_read;                                                        // ddr2_bot_s1_translator:av_read -> ddr2_bot:local_read_req
	wire   [63:0] ddr2_bot_s1_translator_avalon_anti_slave_0_readdata;                                                    // ddr2_bot:local_rdata -> ddr2_bot_s1_translator:av_readdata
	wire          ddr2_bot_s1_translator_avalon_anti_slave_0_readdatavalid;                                               // ddr2_bot:local_rdata_valid -> ddr2_bot_s1_translator:av_readdatavalid
	wire    [7:0] ddr2_bot_s1_translator_avalon_anti_slave_0_byteenable;                                                  // ddr2_bot_s1_translator:av_byteenable -> ddr2_bot:local_be
	wire          ddr2_bot_reset_request_n_reset;                                                                         // ddr2_bot:reset_request_n -> [ddr2_bot_s1_translator:reset, ddr2_bot_s1_translator_avalon_universal_slave_0_agent:reset, ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_020:reset, rsp_xbar_demux_020:reset, rst_controller:reset_in4, rst_controller_002:reset_in4, rst_controller_003:reset_in4, rst_controller_004:reset_in4, rst_controller_005:reset_in4, rst_controller_006:reset_in0, width_adapter_014:reset, width_adapter_015:reset]
	wire          fir_dma_write_master_translator_avalon_universal_master_0_waitrequest;                                  // fir_dma_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> fir_dma_write_master_translator:uav_waitrequest
	wire    [4:0] fir_dma_write_master_translator_avalon_universal_master_0_burstcount;                                   // fir_dma_write_master_translator:uav_burstcount -> fir_dma_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] fir_dma_write_master_translator_avalon_universal_master_0_writedata;                                    // fir_dma_write_master_translator:uav_writedata -> fir_dma_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] fir_dma_write_master_translator_avalon_universal_master_0_address;                                      // fir_dma_write_master_translator:uav_address -> fir_dma_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          fir_dma_write_master_translator_avalon_universal_master_0_lock;                                         // fir_dma_write_master_translator:uav_lock -> fir_dma_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          fir_dma_write_master_translator_avalon_universal_master_0_write;                                        // fir_dma_write_master_translator:uav_write -> fir_dma_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          fir_dma_write_master_translator_avalon_universal_master_0_read;                                         // fir_dma_write_master_translator:uav_read -> fir_dma_write_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] fir_dma_write_master_translator_avalon_universal_master_0_readdata;                                     // fir_dma_write_master_translator_avalon_universal_master_0_agent:av_readdata -> fir_dma_write_master_translator:uav_readdata
	wire          fir_dma_write_master_translator_avalon_universal_master_0_debugaccess;                                  // fir_dma_write_master_translator:uav_debugaccess -> fir_dma_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] fir_dma_write_master_translator_avalon_universal_master_0_byteenable;                                   // fir_dma_write_master_translator:uav_byteenable -> fir_dma_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          fir_dma_write_master_translator_avalon_universal_master_0_readdatavalid;                                // fir_dma_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> fir_dma_write_master_translator:uav_readdatavalid
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest;                              // ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> ddr2_top_clock_bridge_m0_translator:uav_waitrequest
	wire    [4:0] ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_burstcount;                               // ddr2_top_clock_bridge_m0_translator:uav_burstcount -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [127:0] ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_writedata;                                // ddr2_top_clock_bridge_m0_translator:uav_writedata -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_address;                                  // ddr2_top_clock_bridge_m0_translator:uav_address -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_lock;                                     // ddr2_top_clock_bridge_m0_translator:uav_lock -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_write;                                    // ddr2_top_clock_bridge_m0_translator:uav_write -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_read;                                     // ddr2_top_clock_bridge_m0_translator:uav_read -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire  [127:0] ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_readdata;                                 // ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> ddr2_top_clock_bridge_m0_translator:uav_readdata
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess;                              // ddr2_top_clock_bridge_m0_translator:uav_debugaccess -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [15:0] ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_byteenable;                               // ddr2_top_clock_bridge_m0_translator:uav_byteenable -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                            // ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> ddr2_top_clock_bridge_m0_translator:uav_readdatavalid
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // ddr2_top_s1_translator:uav_waitrequest -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [5:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_top_s1_translator:uav_burstcount
	wire   [63:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_top_s1_translator:uav_writedata
	wire   [31:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_top_s1_translator:uav_address
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_top_s1_translator:uav_write
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_top_s1_translator:uav_lock
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_top_s1_translator:uav_read
	wire   [63:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // ddr2_top_s1_translator:uav_readdata -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // ddr2_top_s1_translator:uav_readdatavalid -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_top_s1_translator:uav_debugaccess
	wire    [7:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // ddr2_top_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_top_s1_translator:uav_byteenable
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [138:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [138:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [65:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                             // ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [65:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                              // ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                             // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fir_dma_read_master_translator_avalon_universal_master_0_waitrequest;                                   // fir_dma_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> fir_dma_read_master_translator:uav_waitrequest
	wire    [2:0] fir_dma_read_master_translator_avalon_universal_master_0_burstcount;                                    // fir_dma_read_master_translator:uav_burstcount -> fir_dma_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] fir_dma_read_master_translator_avalon_universal_master_0_writedata;                                     // fir_dma_read_master_translator:uav_writedata -> fir_dma_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] fir_dma_read_master_translator_avalon_universal_master_0_address;                                       // fir_dma_read_master_translator:uav_address -> fir_dma_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          fir_dma_read_master_translator_avalon_universal_master_0_lock;                                          // fir_dma_read_master_translator:uav_lock -> fir_dma_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          fir_dma_read_master_translator_avalon_universal_master_0_write;                                         // fir_dma_read_master_translator:uav_write -> fir_dma_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          fir_dma_read_master_translator_avalon_universal_master_0_read;                                          // fir_dma_read_master_translator:uav_read -> fir_dma_read_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] fir_dma_read_master_translator_avalon_universal_master_0_readdata;                                      // fir_dma_read_master_translator_avalon_universal_master_0_agent:av_readdata -> fir_dma_read_master_translator:uav_readdata
	wire          fir_dma_read_master_translator_avalon_universal_master_0_debugaccess;                                   // fir_dma_read_master_translator:uav_debugaccess -> fir_dma_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] fir_dma_read_master_translator_avalon_universal_master_0_byteenable;                                    // fir_dma_read_master_translator:uav_byteenable -> fir_dma_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          fir_dma_read_master_translator_avalon_universal_master_0_readdatavalid;                                 // fir_dma_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> fir_dma_read_master_translator:uav_readdatavalid
	wire          cpu_data_master_translator_avalon_universal_master_0_waitrequest;                                       // cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	wire    [2:0] cpu_data_master_translator_avalon_universal_master_0_burstcount;                                        // cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_writedata;                                         // cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_address;                                           // cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_data_master_translator_avalon_universal_master_0_lock;                                              // cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_data_master_translator_avalon_universal_master_0_write;                                             // cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_data_master_translator_avalon_universal_master_0_read;                                              // cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_data_master_translator_avalon_universal_master_0_readdata;                                          // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	wire          cpu_data_master_translator_avalon_universal_master_0_debugaccess;                                       // cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_data_master_translator_avalon_universal_master_0_byteenable;                                        // cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_data_master_translator_avalon_universal_master_0_readdatavalid;                                     // cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_waitrequest;                                // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	wire    [2:0] cpu_instruction_master_translator_avalon_universal_master_0_burstcount;                                 // cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_writedata;                                  // cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_address;                                    // cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire          cpu_instruction_master_translator_avalon_universal_master_0_lock;                                       // cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire          cpu_instruction_master_translator_avalon_universal_master_0_write;                                      // cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire          cpu_instruction_master_translator_avalon_universal_master_0_read;                                       // cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] cpu_instruction_master_translator_avalon_universal_master_0_readdata;                                   // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	wire          cpu_instruction_master_translator_avalon_universal_master_0_debugaccess;                                // cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] cpu_instruction_master_translator_avalon_universal_master_0_byteenable;                                 // cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid;                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	wire          dma_0_read_master_translator_avalon_universal_master_0_waitrequest;                                     // dma_0_read_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_0_read_master_translator:uav_waitrequest
	wire    [4:0] dma_0_read_master_translator_avalon_universal_master_0_burstcount;                                      // dma_0_read_master_translator:uav_burstcount -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [127:0] dma_0_read_master_translator_avalon_universal_master_0_writedata;                                       // dma_0_read_master_translator:uav_writedata -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dma_0_read_master_translator_avalon_universal_master_0_address;                                         // dma_0_read_master_translator:uav_address -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_0_read_master_translator_avalon_universal_master_0_lock;                                            // dma_0_read_master_translator:uav_lock -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_0_read_master_translator_avalon_universal_master_0_write;                                           // dma_0_read_master_translator:uav_write -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_0_read_master_translator_avalon_universal_master_0_read;                                            // dma_0_read_master_translator:uav_read -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_read
	wire  [127:0] dma_0_read_master_translator_avalon_universal_master_0_readdata;                                        // dma_0_read_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_0_read_master_translator:uav_readdata
	wire          dma_0_read_master_translator_avalon_universal_master_0_debugaccess;                                     // dma_0_read_master_translator:uav_debugaccess -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [15:0] dma_0_read_master_translator_avalon_universal_master_0_byteenable;                                      // dma_0_read_master_translator:uav_byteenable -> dma_0_read_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_0_read_master_translator_avalon_universal_master_0_readdatavalid;                                   // dma_0_read_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_0_read_master_translator:uav_readdatavalid
	wire          dma_0_write_master_translator_avalon_universal_master_0_waitrequest;                                    // dma_0_write_master_translator_avalon_universal_master_0_agent:av_waitrequest -> dma_0_write_master_translator:uav_waitrequest
	wire    [4:0] dma_0_write_master_translator_avalon_universal_master_0_burstcount;                                     // dma_0_write_master_translator:uav_burstcount -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [127:0] dma_0_write_master_translator_avalon_universal_master_0_writedata;                                      // dma_0_write_master_translator:uav_writedata -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] dma_0_write_master_translator_avalon_universal_master_0_address;                                        // dma_0_write_master_translator:uav_address -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_address
	wire          dma_0_write_master_translator_avalon_universal_master_0_lock;                                           // dma_0_write_master_translator:uav_lock -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_lock
	wire          dma_0_write_master_translator_avalon_universal_master_0_write;                                          // dma_0_write_master_translator:uav_write -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_write
	wire          dma_0_write_master_translator_avalon_universal_master_0_read;                                           // dma_0_write_master_translator:uav_read -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_read
	wire  [127:0] dma_0_write_master_translator_avalon_universal_master_0_readdata;                                       // dma_0_write_master_translator_avalon_universal_master_0_agent:av_readdata -> dma_0_write_master_translator:uav_readdata
	wire          dma_0_write_master_translator_avalon_universal_master_0_debugaccess;                                    // dma_0_write_master_translator:uav_debugaccess -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [15:0] dma_0_write_master_translator_avalon_universal_master_0_byteenable;                                     // dma_0_write_master_translator:uav_byteenable -> dma_0_write_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          dma_0_write_master_translator_avalon_universal_master_0_readdatavalid;                                  // dma_0_write_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> dma_0_write_master_translator:uav_readdatavalid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // flash_ssram_pipeline_bridge_s0_translator:uav_waitrequest -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> flash_ssram_pipeline_bridge_s0_translator:uav_burstcount
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                  // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> flash_ssram_pipeline_bridge_s0_translator:uav_writedata
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                    // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> flash_ssram_pipeline_bridge_s0_translator:uav_address
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                      // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> flash_ssram_pipeline_bridge_s0_translator:uav_write
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                       // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> flash_ssram_pipeline_bridge_s0_translator:uav_lock
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                       // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> flash_ssram_pipeline_bridge_s0_translator:uav_read
	wire   [31:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                   // flash_ssram_pipeline_bridge_s0_translator:uav_readdata -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // flash_ssram_pipeline_bridge_s0_translator:uav_readdatavalid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> flash_ssram_pipeline_bridge_s0_translator:uav_debugaccess
	wire    [3:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> flash_ssram_pipeline_bridge_s0_translator:uav_byteenable
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;               // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;               // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;          // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;           // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;          // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // slow_peripheral_bridge_s0_translator:uav_waitrequest -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> slow_peripheral_bridge_s0_translator:uav_burstcount
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                       // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> slow_peripheral_bridge_s0_translator:uav_writedata
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                         // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> slow_peripheral_bridge_s0_translator:uav_address
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> slow_peripheral_bridge_s0_translator:uav_write
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> slow_peripheral_bridge_s0_translator:uav_lock
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> slow_peripheral_bridge_s0_translator:uav_read
	wire   [31:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                        // slow_peripheral_bridge_s0_translator:uav_readdata -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // slow_peripheral_bridge_s0_translator:uav_readdatavalid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> slow_peripheral_bridge_s0_translator:uav_debugaccess
	wire    [3:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> slow_peripheral_bridge_s0_translator:uav_byteenable
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                     // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;               // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;               // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // ddr2_top_clock_bridge_s0_translator:uav_waitrequest -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [4:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_top_clock_bridge_s0_translator:uav_burstcount
	wire  [127:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                        // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_top_clock_bridge_s0_translator:uav_writedata
	wire   [31:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                          // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_top_clock_bridge_s0_translator:uav_address
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                            // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_top_clock_bridge_s0_translator:uav_write
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                             // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_top_clock_bridge_s0_translator:uav_lock
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                             // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_top_clock_bridge_s0_translator:uav_read
	wire  [127:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                         // ddr2_top_clock_bridge_s0_translator:uav_readdata -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // ddr2_top_clock_bridge_s0_translator:uav_readdatavalid -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_top_clock_bridge_s0_translator:uav_debugaccess
	wire   [15:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_top_clock_bridge_s0_translator:uav_byteenable
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [215:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                      // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [215:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [129:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [129:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // cpu_jtag_debug_module_translator:uav_waitrequest -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_jtag_debug_module_translator:uav_burstcount
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;                           // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_jtag_debug_module_translator:uav_writedata
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_jtag_debug_module_translator:uav_address
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_jtag_debug_module_translator:uav_write
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_jtag_debug_module_translator:uav_lock
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_jtag_debug_module_translator:uav_read
	wire   [31:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                            // cpu_jtag_debug_module_translator:uav_readdata -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // cpu_jtag_debug_module_translator:uav_readdatavalid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_jtag_debug_module_translator:uav_debugaccess
	wire    [3:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_jtag_debug_module_translator:uav_byteenable
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                    // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                   // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // ddr2_bot_clock_bridge_s0_translator:uav_waitrequest -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [4:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_bot_clock_bridge_s0_translator:uav_burstcount
	wire  [127:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata;                        // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_bot_clock_bridge_s0_translator:uav_writedata
	wire   [31:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address;                          // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_bot_clock_bridge_s0_translator:uav_address
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write;                            // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_bot_clock_bridge_s0_translator:uav_write
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock;                             // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_bot_clock_bridge_s0_translator:uav_lock
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read;                             // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_bot_clock_bridge_s0_translator:uav_read
	wire  [127:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata;                         // ddr2_bot_clock_bridge_s0_translator:uav_readdata -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // ddr2_bot_clock_bridge_s0_translator:uav_readdatavalid -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_bot_clock_bridge_s0_translator:uav_debugaccess
	wire   [15:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_bot_clock_bridge_s0_translator:uav_byteenable
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [215:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data;                      // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [215:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire  [129:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [129:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // dma_0_control_port_slave_translator:uav_waitrequest -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> dma_0_control_port_slave_translator:uav_burstcount
	wire   [31:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                        // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> dma_0_control_port_slave_translator:uav_writedata
	wire   [31:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address;                          // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_address -> dma_0_control_port_slave_translator:uav_address
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write;                            // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_write -> dma_0_control_port_slave_translator:uav_write
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock;                             // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_lock -> dma_0_control_port_slave_translator:uav_lock
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read;                             // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_read -> dma_0_control_port_slave_translator:uav_read
	wire   [31:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                         // dma_0_control_port_slave_translator:uav_readdata -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // dma_0_control_port_slave_translator:uav_readdatavalid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dma_0_control_port_slave_translator:uav_debugaccess
	wire    [3:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> dma_0_control_port_slave_translator:uav_byteenable
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [107:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                      // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [107:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest;                             // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> slow_peripheral_bridge_m0_translator:uav_waitrequest
	wire    [2:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount;                              // slow_peripheral_bridge_m0_translator:uav_burstcount -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata;                               // slow_peripheral_bridge_m0_translator:uav_writedata -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire    [9:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address;                                 // slow_peripheral_bridge_m0_translator:uav_address -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock;                                    // slow_peripheral_bridge_m0_translator:uav_lock -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write;                                   // slow_peripheral_bridge_m0_translator:uav_write -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read;                                    // slow_peripheral_bridge_m0_translator:uav_read -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata;                                // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> slow_peripheral_bridge_m0_translator:uav_readdata
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess;                             // slow_peripheral_bridge_m0_translator:uav_debugaccess -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable;                              // slow_peripheral_bridge_m0_translator:uav_byteenable -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                           // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> slow_peripheral_bridge_m0_translator:uav_readdatavalid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                             // high_res_timer_s1_translator:uav_waitrequest -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                              // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> high_res_timer_s1_translator:uav_burstcount
	wire   [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                               // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> high_res_timer_s1_translator:uav_writedata
	wire    [9:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                 // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> high_res_timer_s1_translator:uav_address
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> high_res_timer_s1_translator:uav_write
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> high_res_timer_s1_translator:uav_lock
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> high_res_timer_s1_translator:uav_read
	wire   [31:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                // high_res_timer_s1_translator:uav_readdata -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                           // high_res_timer_s1_translator:uav_readdatavalid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                             // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> high_res_timer_s1_translator:uav_debugaccess
	wire    [3:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                              // high_res_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> high_res_timer_s1_translator:uav_byteenable
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                      // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                             // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                            // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                         // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                 // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                          // high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                         // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                       // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                        // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                       // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                   // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire    [9:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                      // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                 // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // performance_counter_control_slave_translator:uav_waitrequest -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;              // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> performance_counter_control_slave_translator:uav_burstcount
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;               // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> performance_counter_control_slave_translator:uav_writedata
	wire    [9:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                 // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> performance_counter_control_slave_translator:uav_address
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                   // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> performance_counter_control_slave_translator:uav_write
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> performance_counter_control_slave_translator:uav_lock
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> performance_counter_control_slave_translator:uav_read
	wire   [31:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                // performance_counter_control_slave_translator:uav_readdata -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // performance_counter_control_slave_translator:uav_readdatavalid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> performance_counter_control_slave_translator:uav_debugaccess
	wire    [3:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;              // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> performance_counter_control_slave_translator:uav_byteenable
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;             // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;            // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // sys_clk_timer_s1_translator:uav_waitrequest -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sys_clk_timer_s1_translator:uav_burstcount
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sys_clk_timer_s1_translator:uav_writedata
	wire    [9:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_address -> sys_clk_timer_s1_translator:uav_address
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_write -> sys_clk_timer_s1_translator:uav_write
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sys_clk_timer_s1_translator:uav_lock
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_read -> sys_clk_timer_s1_translator:uav_read
	wire   [31:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // sys_clk_timer_s1_translator:uav_readdata -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // sys_clk_timer_s1_translator:uav_readdatavalid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sys_clk_timer_s1_translator:uav_debugaccess
	wire    [3:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sys_clk_timer_s1_translator:uav_byteenable
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // sysid_control_slave_translator:uav_waitrequest -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_control_slave_translator:uav_burstcount
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                             // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_control_slave_translator:uav_writedata
	wire    [9:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                               // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_control_slave_translator:uav_address
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_control_slave_translator:uav_write
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_control_slave_translator:uav_lock
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_control_slave_translator:uav_read
	wire   [31:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                              // sysid_control_slave_translator:uav_readdata -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // sysid_control_slave_translator:uav_readdatavalid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_control_slave_translator:uav_debugaccess
	wire    [3:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // sysid_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_control_slave_translator:uav_byteenable
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // sysid_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // fir_dma_control_translator:uav_waitrequest -> fir_dma_control_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] fir_dma_control_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // fir_dma_control_translator_avalon_universal_slave_0_agent:m0_burstcount -> fir_dma_control_translator:uav_burstcount
	wire   [31:0] fir_dma_control_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // fir_dma_control_translator_avalon_universal_slave_0_agent:m0_writedata -> fir_dma_control_translator:uav_writedata
	wire    [9:0] fir_dma_control_translator_avalon_universal_slave_0_agent_m0_address;                                   // fir_dma_control_translator_avalon_universal_slave_0_agent:m0_address -> fir_dma_control_translator:uav_address
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_m0_write;                                     // fir_dma_control_translator_avalon_universal_slave_0_agent:m0_write -> fir_dma_control_translator:uav_write
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_m0_lock;                                      // fir_dma_control_translator_avalon_universal_slave_0_agent:m0_lock -> fir_dma_control_translator:uav_lock
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_m0_read;                                      // fir_dma_control_translator_avalon_universal_slave_0_agent:m0_read -> fir_dma_control_translator:uav_read
	wire   [31:0] fir_dma_control_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // fir_dma_control_translator:uav_readdata -> fir_dma_control_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // fir_dma_control_translator:uav_readdatavalid -> fir_dma_control_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // fir_dma_control_translator_avalon_universal_slave_0_agent:m0_debugaccess -> fir_dma_control_translator:uav_debugaccess
	wire    [3:0] fir_dma_control_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // fir_dma_control_translator_avalon_universal_slave_0_agent:m0_byteenable -> fir_dma_control_translator:uav_byteenable
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // fir_dma_control_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // fir_dma_control_translator_avalon_universal_slave_0_agent:rf_source_valid -> fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // fir_dma_control_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_data;                               // fir_dma_control_translator_avalon_universal_slave_0_agent:rf_source_data -> fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> fir_dma_control_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> fir_dma_control_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> fir_dma_control_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> fir_dma_control_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> fir_dma_control_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // fir_dma_control_translator_avalon_universal_slave_0_agent:rf_sink_ready -> fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // fir_dma_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // fir_dma_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> fir_dma_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                         // fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> fir_dma_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                          // fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> fir_dma_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                         // fir_dma_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // pll_pll_slave_translator:uav_waitrequest -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> pll_pll_slave_translator:uav_burstcount
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> pll_pll_slave_translator:uav_writedata
	wire    [9:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address;                                     // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_address -> pll_pll_slave_translator:uav_address
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write;                                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_write -> pll_pll_slave_translator:uav_write
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock;                                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_lock -> pll_pll_slave_translator:uav_lock
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read;                                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_read -> pll_pll_slave_translator:uav_read
	wire   [31:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // pll_pll_slave_translator:uav_readdata -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // pll_pll_slave_translator:uav_readdatavalid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pll_pll_slave_translator:uav_debugaccess
	wire    [3:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // pll_pll_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> pll_pll_slave_translator:uav_byteenable
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // pll_pll_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                            // pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                           // pll_pll_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // button_pio_s1_translator:uav_waitrequest -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_pio_s1_translator:uav_burstcount
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_pio_s1_translator:uav_writedata
	wire    [9:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_pio_s1_translator:uav_address
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_pio_s1_translator:uav_write
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_pio_s1_translator:uav_lock
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_pio_s1_translator:uav_read
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // button_pio_s1_translator:uav_readdata -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // button_pio_s1_translator:uav_readdatavalid -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_pio_s1_translator:uav_debugaccess
	wire    [3:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_pio_s1_translator:uav_byteenable
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                    // led_pio_s1_translator:uav_waitrequest -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_pio_s1_translator:uav_burstcount
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                      // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_pio_s1_translator:uav_writedata
	wire    [9:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                        // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_pio_s1_translator:uav_address
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                          // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_pio_s1_translator:uav_write
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                           // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_pio_s1_translator:uav_lock
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                           // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_pio_s1_translator:uav_read
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                       // led_pio_s1_translator:uav_readdata -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                  // led_pio_s1_translator:uav_readdatavalid -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_pio_s1_translator:uav_debugaccess
	wire    [3:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_pio_s1_translator:uav_byteenable
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                             // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                   // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                           // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                   // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                          // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                        // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                 // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                              // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                               // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                              // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // lcd_display_control_slave_translator:uav_waitrequest -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_display_control_slave_translator:uav_burstcount
	wire   [31:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                       // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_display_control_slave_translator:uav_writedata
	wire    [9:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                         // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_display_control_slave_translator:uav_address
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                           // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_display_control_slave_translator:uav_write
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                            // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_display_control_slave_translator:uav_lock
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                            // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_display_control_slave_translator:uav_read
	wire   [31:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                        // lcd_display_control_slave_translator:uav_readdata -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // lcd_display_control_slave_translator:uav_readdatavalid -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_display_control_slave_translator:uav_debugaccess
	wire    [3:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_display_control_slave_translator:uav_byteenable
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                     // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // seven_seg_pio_s1_translator:uav_waitrequest -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> seven_seg_pio_s1_translator:uav_burstcount
	wire   [31:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> seven_seg_pio_s1_translator:uav_writedata
	wire    [9:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> seven_seg_pio_s1_translator:uav_address
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> seven_seg_pio_s1_translator:uav_write
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> seven_seg_pio_s1_translator:uav_lock
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> seven_seg_pio_s1_translator:uav_read
	wire   [31:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // seven_seg_pio_s1_translator:uav_readdata -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // seven_seg_pio_s1_translator:uav_readdatavalid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> seven_seg_pio_s1_translator:uav_debugaccess
	wire    [3:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> seven_seg_pio_s1_translator:uav_byteenable
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [83:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [83:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_waitrequest;                        // flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> flash_ssram_pipeline_bridge_m0_translator:uav_waitrequest
	wire    [2:0] flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_burstcount;                         // flash_ssram_pipeline_bridge_m0_translator:uav_burstcount -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_writedata;                          // flash_ssram_pipeline_bridge_m0_translator:uav_writedata -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [26:0] flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_address;                            // flash_ssram_pipeline_bridge_m0_translator:uav_address -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_lock;                               // flash_ssram_pipeline_bridge_m0_translator:uav_lock -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_write;                              // flash_ssram_pipeline_bridge_m0_translator:uav_write -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_read;                               // flash_ssram_pipeline_bridge_m0_translator:uav_read -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_readdata;                           // flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> flash_ssram_pipeline_bridge_m0_translator:uav_readdata
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_debugaccess;                        // flash_ssram_pipeline_bridge_m0_translator:uav_debugaccess -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_byteenable;                         // flash_ssram_pipeline_bridge_m0_translator:uav_byteenable -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                      // flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> flash_ssram_pipeline_bridge_m0_translator:uav_readdatavalid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                     // ssram_uas_translator:uav_waitrequest -> ssram_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                      // ssram_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> ssram_uas_translator:uav_burstcount
	wire   [31:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                       // ssram_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> ssram_uas_translator:uav_writedata
	wire   [26:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_address;                                         // ssram_uas_translator_avalon_universal_slave_0_agent:m0_address -> ssram_uas_translator:uav_address
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_write;                                           // ssram_uas_translator_avalon_universal_slave_0_agent:m0_write -> ssram_uas_translator:uav_write
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                            // ssram_uas_translator_avalon_universal_slave_0_agent:m0_lock -> ssram_uas_translator:uav_lock
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_read;                                            // ssram_uas_translator_avalon_universal_slave_0_agent:m0_read -> ssram_uas_translator:uav_read
	wire   [31:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                        // ssram_uas_translator:uav_readdata -> ssram_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                   // ssram_uas_translator:uav_readdatavalid -> ssram_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                     // ssram_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ssram_uas_translator:uav_debugaccess
	wire    [3:0] ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                      // ssram_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> ssram_uas_translator:uav_byteenable
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                              // ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                                    // ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                            // ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [94:0] ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                     // ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                                    // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                           // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                                 // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                         // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [94:0] ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                  // ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                                 // ssram_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                               // ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                                // ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                               // ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ssram_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // ext_flash_uas_translator:uav_waitrequest -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> ext_flash_uas_translator:uav_burstcount
	wire   [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> ext_flash_uas_translator:uav_writedata
	wire   [26:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address;                                     // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_address -> ext_flash_uas_translator:uav_address
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write;                                       // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_write -> ext_flash_uas_translator:uav_write
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock;                                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_lock -> ext_flash_uas_translator:uav_lock
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read;                                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_read -> ext_flash_uas_translator:uav_read
	wire   [15:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // ext_flash_uas_translator:uav_readdata -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // ext_flash_uas_translator:uav_readdatavalid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ext_flash_uas_translator:uav_debugaccess
	wire    [1:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // ext_flash_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> ext_flash_uas_translator:uav_byteenable
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire   [76:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire   [76:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // ext_flash_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                           // ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                            // ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                           // ext_flash_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest;                              // ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_waitrequest -> ddr2_bot_clock_bridge_m0_translator:uav_waitrequest
	wire    [4:0] ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_burstcount;                               // ddr2_bot_clock_bridge_m0_translator:uav_burstcount -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [127:0] ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_writedata;                                // ddr2_bot_clock_bridge_m0_translator:uav_writedata -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [26:0] ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_address;                                  // ddr2_bot_clock_bridge_m0_translator:uav_address -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_address
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_lock;                                     // ddr2_bot_clock_bridge_m0_translator:uav_lock -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_lock
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_write;                                    // ddr2_bot_clock_bridge_m0_translator:uav_write -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_write
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_read;                                     // ddr2_bot_clock_bridge_m0_translator:uav_read -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_read
	wire  [127:0] ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_readdata;                                 // ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdata -> ddr2_bot_clock_bridge_m0_translator:uav_readdata
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess;                              // ddr2_bot_clock_bridge_m0_translator:uav_debugaccess -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [15:0] ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_byteenable;                               // ddr2_bot_clock_bridge_m0_translator:uav_byteenable -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid;                            // ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:av_readdatavalid -> ddr2_bot_clock_bridge_m0_translator:uav_readdatavalid
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // ddr2_bot_s1_translator:uav_waitrequest -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [5:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> ddr2_bot_s1_translator:uav_burstcount
	wire   [63:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> ddr2_bot_s1_translator:uav_writedata
	wire   [26:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_address -> ddr2_bot_s1_translator:uav_address
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_write -> ddr2_bot_s1_translator:uav_write
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_lock -> ddr2_bot_s1_translator:uav_lock
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_read -> ddr2_bot_s1_translator:uav_read
	wire   [63:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // ddr2_bot_s1_translator:uav_readdata -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // ddr2_bot_s1_translator:uav_readdatavalid -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ddr2_bot_s1_translator:uav_debugaccess
	wire    [7:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> ddr2_bot_s1_translator:uav_byteenable
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [133:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [133:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [65:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                             // ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [65:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                              // ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                             // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                         // fir_dma_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_valid;                               // fir_dma_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                       // fir_dma_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [101:0] fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_data;                                // fir_dma_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_ready;                               // addr_router:sink_ready -> fir_dma_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                     // ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                           // ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                   // ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [209:0] ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                            // ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire          ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                           // addr_router_001:sink_ready -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [137:0] ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // ddr2_top_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router:sink_ready -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                          // fir_dma_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_valid;                                // fir_dma_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_002:sink_valid
	wire          fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                        // fir_dma_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [106:0] fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_data;                                 // fir_dma_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_002:sink_data
	wire          fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_ready;                                // addr_router_002:sink_ready -> fir_dma_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                              // cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid;                                    // cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_003:sink_valid
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                            // cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [106:0] cpu_data_master_translator_avalon_universal_master_0_agent_cp_data;                                     // cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_003:sink_data
	wire          cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready;                                    // addr_router_003:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                       // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                             // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_004:sink_valid
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                     // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [106:0] cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_004:sink_data
	wire          cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                             // addr_router_004:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                            // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid;                                  // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                          // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [214:0] dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data;                                   // dma_0_read_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready;                                  // addr_router_005:sink_ready -> dma_0_read_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                           // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_006:sink_endofpacket
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid;                                 // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_006:sink_valid
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                         // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_006:sink_startofpacket
	wire  [214:0] dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data;                                  // dma_0_write_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_006:sink_data
	wire          dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready;                                 // addr_router_006:sink_ready -> dma_0_write_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                      // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [106:0] flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                       // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_001:sink_ready -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                           // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [106:0] slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                            // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_002:sink_ready -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                            // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [214:0] ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                             // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_003:sink_ready -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                               // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [106:0] cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                                // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_004:sink_ready -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid;                            // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [214:0] ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data;                             // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_005:sink_ready -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid;                            // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [106:0] dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data;                             // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_006:sink_ready -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                    // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_007:sink_endofpacket
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                          // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_007:sink_valid
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                  // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_007:sink_startofpacket
	wire   [82:0] slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                           // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_007:sink_data
	wire          slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                          // addr_router_007:sink_ready -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                             // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                   // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                           // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire   [82:0] high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                    // high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                   // id_router_007:sink_ready -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                   // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire   [82:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                         // id_router_008:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                   // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire   [82:0] performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                    // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_009:sink_ready -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire   [82:0] sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_010:sink_ready -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                 // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire   [82:0] sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                                  // sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire          sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_011:sink_ready -> sysid_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // fir_dma_control_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rp_valid;                                     // fir_dma_control_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // fir_dma_control_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire   [82:0] fir_dma_control_translator_avalon_universal_slave_0_agent_rp_data;                                      // fir_dma_control_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire          fir_dma_control_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_012:sink_ready -> fir_dma_control_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid;                                       // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire   [82:0] pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data;                                        // pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire          pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_013:sink_ready -> pll_pll_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	wire   [82:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_014:sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                    // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                          // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                  // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	wire   [82:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                           // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                          // id_router_015:sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                           // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	wire   [82:0] lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                            // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	wire          lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_016:sink_ready -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	wire   [82:0] seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	wire          seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_017:sink_ready -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;               // flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_008:sink_endofpacket
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                     // flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_008:sink_valid
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;             // flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_008:sink_startofpacket
	wire   [93:0] flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                      // flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_008:sink_data
	wire          flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router_008:sink_ready -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                     // ssram_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                           // ssram_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                   // ssram_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	wire   [93:0] ssram_uas_translator_avalon_universal_slave_0_agent_rp_data;                                            // ssram_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	wire          ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                           // id_router_018:sink_ready -> ssram_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid;                                       // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	wire   [75:0] ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data;                                        // ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	wire          ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_019:sink_ready -> ext_flash_uas_translator_avalon_universal_slave_0_agent:rp_ready
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket;                     // ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_009:sink_endofpacket
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid;                           // ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_009:sink_valid
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket;                   // ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_009:sink_startofpacket
	wire  [204:0] ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data;                            // ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_data -> addr_router_009:sink_data
	wire          ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready;                           // addr_router_009:sink_ready -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:cp_ready
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	wire  [132:0] ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	wire          ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_020:sink_ready -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_003_src_endofpacket;                                                                        // addr_router_003:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_003_src_valid;                                                                              // addr_router_003:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_003_src_startofpacket;                                                                      // addr_router_003:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [106:0] addr_router_003_src_data;                                                                               // addr_router_003:src_data -> limiter:cmd_sink_data
	wire    [5:0] addr_router_003_src_channel;                                                                            // addr_router_003:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_003_src_ready;                                                                              // limiter:cmd_sink_ready -> addr_router_003:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                            // limiter:rsp_src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                                  // limiter:rsp_src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                          // limiter:rsp_src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_rsp_src_data;                                                                                   // limiter:rsp_src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_rsp_src_channel;                                                                                // limiter:rsp_src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                                  // cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_004_src_endofpacket;                                                                        // addr_router_004:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_004_src_valid;                                                                              // addr_router_004:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_004_src_startofpacket;                                                                      // addr_router_004:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [106:0] addr_router_004_src_data;                                                                               // addr_router_004:src_data -> limiter_001:cmd_sink_data
	wire    [5:0] addr_router_004_src_channel;                                                                            // addr_router_004:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_004_src_ready;                                                                              // limiter_001:cmd_sink_ready -> addr_router_004:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                        // limiter_001:rsp_src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                              // limiter_001:rsp_src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                      // limiter_001:rsp_src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] limiter_001_rsp_src_data;                                                                               // limiter_001:rsp_src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] limiter_001_rsp_src_channel;                                                                            // limiter_001:rsp_src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_001_rsp_src_ready;                                                                              // cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_007_src_endofpacket;                                                                        // addr_router_007:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_007_src_valid;                                                                              // addr_router_007:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_007_src_startofpacket;                                                                      // addr_router_007:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire   [82:0] addr_router_007_src_data;                                                                               // addr_router_007:src_data -> limiter_002:cmd_sink_data
	wire   [10:0] addr_router_007_src_channel;                                                                            // addr_router_007:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_007_src_ready;                                                                              // limiter_002:cmd_sink_ready -> addr_router_007:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                        // limiter_002:rsp_src_endofpacket -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                              // limiter_002:rsp_src_valid -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                      // limiter_002:rsp_src_startofpacket -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [82:0] limiter_002_rsp_src_data;                                                                               // limiter_002:rsp_src_data -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire   [10:0] limiter_002_rsp_src_channel;                                                                            // limiter_002:rsp_src_channel -> slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_002_rsp_src_ready;                                                                              // slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_002:rsp_src_ready
	wire          addr_router_008_src_endofpacket;                                                                        // addr_router_008:src_endofpacket -> limiter_003:cmd_sink_endofpacket
	wire          addr_router_008_src_valid;                                                                              // addr_router_008:src_valid -> limiter_003:cmd_sink_valid
	wire          addr_router_008_src_startofpacket;                                                                      // addr_router_008:src_startofpacket -> limiter_003:cmd_sink_startofpacket
	wire   [93:0] addr_router_008_src_data;                                                                               // addr_router_008:src_data -> limiter_003:cmd_sink_data
	wire    [1:0] addr_router_008_src_channel;                                                                            // addr_router_008:src_channel -> limiter_003:cmd_sink_channel
	wire          addr_router_008_src_ready;                                                                              // limiter_003:cmd_sink_ready -> addr_router_008:src_ready
	wire          limiter_003_rsp_src_endofpacket;                                                                        // limiter_003:rsp_src_endofpacket -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_003_rsp_src_valid;                                                                              // limiter_003:rsp_src_valid -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_003_rsp_src_startofpacket;                                                                      // limiter_003:rsp_src_startofpacket -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire   [93:0] limiter_003_rsp_src_data;                                                                               // limiter_003:rsp_src_data -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] limiter_003_rsp_src_channel;                                                                            // limiter_003:rsp_src_channel -> flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_003_rsp_src_ready;                                                                              // flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> limiter_003:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                      // burst_adapter:source0_endofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                            // burst_adapter:source0_valid -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                    // burst_adapter:source0_startofpacket -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [75:0] burst_adapter_source0_data;                                                                             // burst_adapter:source0_data -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                            // ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [1:0] burst_adapter_source0_channel;                                                                          // burst_adapter:source0_channel -> ext_flash_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                                         // rst_controller:reset_out -> [ddr2_bot:soft_reset_n, ddr2_top:soft_reset_n]
	wire          cpu_jtag_debug_module_reset_reset;                                                                      // cpu:jtag_debug_module_resetrequest -> [rst_controller:reset_in3, rst_controller_001:reset_in0, rst_controller_002:reset_in3, rst_controller_003:reset_in3, rst_controller_004:reset_in3, rst_controller_005:reset_in3, rst_controller_006:reset_in4]
	wire          rst_controller_001_reset_out_reset;                                                                     // rst_controller_001:reset_out -> [ddr2_bot:global_reset_n, ddr2_top:global_reset_n]
	wire          rst_controller_002_reset_out_reset;                                                                     // rst_controller_002:reset_out -> [addr_router_007:reset, button_pio:reset_n, button_pio_s1_translator:reset, button_pio_s1_translator_avalon_universal_slave_0_agent:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux_007:reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:out_reset, crosser_007:out_reset, high_res_timer:reset_n, high_res_timer_s1_translator:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent:reset, high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, irq_synchronizer_004:receiver_reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_display:reset_n, lcd_display_control_slave_translator:reset, lcd_display_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_pio:reset_n, led_pio_s1_translator:reset, led_pio_s1_translator_avalon_universal_slave_0_agent:reset, led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter_002:reset, performance_counter:reset_n, performance_counter_control_slave_translator:reset, performance_counter_control_slave_translator_avalon_universal_slave_0_agent:reset, performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_mux_007:reset, seven_seg_pio:reset_n, seven_seg_pio_s1_translator:reset, seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:reset, seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, slow_peripheral_bridge:m0_reset, slow_peripheral_bridge_m0_translator:reset, slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent:reset, sys_clk_timer:reset_n, sys_clk_timer_s1_translator:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:reset, sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid:reset_n, sysid_control_slave_translator:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire          rst_controller_003_reset_out_reset;                                                                     // rst_controller_003:reset_out -> [addr_router:reset, addr_router_002:reset, cmd_xbar_demux:reset, cmd_xbar_demux_002:reset, crosser:in_reset, crosser_001:out_reset, crosser_002:in_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_005:out_reset, crosser_006:in_reset, crosser_007:in_reset, fir_dma:reset, fir_dma_control_translator:reset, fir_dma_control_translator_avalon_universal_slave_0_agent:reset, fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, fir_dma_read_master_translator:reset, fir_dma_read_master_translator_avalon_universal_master_0_agent:reset, fir_dma_write_master_translator:reset, fir_dma_write_master_translator_avalon_universal_master_0_agent:reset, id_router_012:reset, id_router_013:reset, irq_synchronizer_003:receiver_reset, pll:reset, pll_pll_slave_translator:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, width_adapter:reset, width_adapter_001:reset]
	wire          rst_controller_004_reset_out_reset;                                                                     // rst_controller_004:reset_out -> [addr_router_003:reset, addr_router_004:reset, addr_router_005:reset, addr_router_006:reset, addr_router_008:reset, burst_adapter:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, cmd_xbar_demux_005:reset, cmd_xbar_demux_006:reset, cmd_xbar_demux_008:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cpu:reset_n, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_jtag_debug_module_translator:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, crosser_002:out_reset, crosser_003:in_reset, ddr2_bot_clock_bridge:s0_reset, ddr2_bot_clock_bridge_s0_translator:reset, ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:reset, ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ddr2_top_clock_bridge:s0_reset, ddr2_top_clock_bridge_s0_translator:reset, ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:reset, ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_0:system_reset_n, dma_0_control_port_slave_translator:reset, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:reset, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, dma_0_read_master_translator:reset, dma_0_read_master_translator_avalon_universal_master_0_agent:reset, dma_0_write_master_translator:reset, dma_0_write_master_translator_avalon_universal_master_0_agent:reset, ext_flash:reset_reset, ext_flash_uas_translator:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, flash_ssram_pipeline_bridge:reset, flash_ssram_pipeline_bridge_m0_translator:reset, flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent:reset, flash_ssram_pipeline_bridge_s0_translator:reset, flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:reset, flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, flash_ssram_tristate_bridge_bridge_0:reset, flash_ssram_tristate_bridge_pinSharer_0:reset_reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_018:reset, id_router_019:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, irq_synchronizer_004:sender_reset, limiter:reset, limiter_001:reset, limiter_003:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_018:reset, rsp_xbar_demux_019:reset, rsp_xbar_mux_003:reset, rsp_xbar_mux_004:reset, rsp_xbar_mux_008:reset, slow_peripheral_bridge:s0_reset, slow_peripheral_bridge_s0_translator:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ssram:reset_reset, ssram_uas_translator:reset, ssram_uas_translator_avalon_universal_slave_0_agent:reset, ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_004:reset, width_adapter_005:reset, width_adapter_006:reset, width_adapter_007:reset, width_adapter_008:reset, width_adapter_009:reset, width_adapter_010:reset, width_adapter_011:reset, width_adapter_012:reset, width_adapter_013:reset]
	wire          rst_controller_005_reset_out_reset;                                                                     // rst_controller_005:reset_out -> [addr_router_001:reset, cmd_xbar_demux_001:reset, ddr2_top_clock_bridge:m0_reset, ddr2_top_clock_bridge_m0_translator:reset, ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_006_reset_out_reset;                                                                     // rst_controller_006:reset_out -> [addr_router_009:reset, cmd_xbar_demux_009:reset, ddr2_bot_clock_bridge:m0_reset, ddr2_bot_clock_bridge_m0_translator:reset, ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:reset]
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                    // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                          // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                                  // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [137:0] cmd_xbar_demux_001_src0_data;                                                                           // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire    [1:0] cmd_xbar_demux_001_src0_channel;                                                                        // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                          // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_src1_endofpacket;                                                                        // rsp_xbar_demux:src1_endofpacket -> width_adapter_003:in_endofpacket
	wire          rsp_xbar_demux_src1_valid;                                                                              // rsp_xbar_demux:src1_valid -> width_adapter_003:in_valid
	wire          rsp_xbar_demux_src1_startofpacket;                                                                      // rsp_xbar_demux:src1_startofpacket -> width_adapter_003:in_startofpacket
	wire  [137:0] rsp_xbar_demux_src1_data;                                                                               // rsp_xbar_demux:src1_data -> width_adapter_003:in_data
	wire    [1:0] rsp_xbar_demux_src1_channel;                                                                            // rsp_xbar_demux:src1_channel -> width_adapter_003:in_channel
	wire          cmd_xbar_mux_src_endofpacket;                                                                           // cmd_xbar_mux:src_endofpacket -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_src_valid;                                                                                 // cmd_xbar_mux:src_valid -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_src_startofpacket;                                                                         // cmd_xbar_mux:src_startofpacket -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [137:0] cmd_xbar_mux_src_data;                                                                                  // cmd_xbar_mux:src_data -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire    [1:0] cmd_xbar_mux_src_channel;                                                                               // cmd_xbar_mux:src_channel -> ddr2_top_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_src_ready;                                                                                 // ddr2_top_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire          id_router_src_endofpacket;                                                                              // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          id_router_src_valid;                                                                                    // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire          id_router_src_startofpacket;                                                                            // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [137:0] id_router_src_data;                                                                                     // id_router:src_data -> rsp_xbar_demux:sink_data
	wire    [1:0] id_router_src_channel;                                                                                  // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire          id_router_src_ready;                                                                                    // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                    // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                          // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_001:sink1_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                                  // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src0_data;                                                                           // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_001:sink1_data
	wire    [5:0] cmd_xbar_demux_003_src0_channel;                                                                        // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_001:sink1_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                          // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_003_src1_endofpacket;                                                                    // cmd_xbar_demux_003:src1_endofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src1_valid;                                                                          // cmd_xbar_demux_003:src1_valid -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src1_startofpacket;                                                                  // cmd_xbar_demux_003:src1_startofpacket -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src1_data;                                                                           // cmd_xbar_demux_003:src1_data -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_demux_003_src1_channel;                                                                        // cmd_xbar_demux_003:src1_channel -> slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_003_src3_endofpacket;                                                                    // cmd_xbar_demux_003:src3_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_003_src3_valid;                                                                          // cmd_xbar_demux_003:src3_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_003_src3_startofpacket;                                                                  // cmd_xbar_demux_003:src3_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src3_data;                                                                           // cmd_xbar_demux_003:src3_data -> cmd_xbar_mux_004:sink0_data
	wire    [5:0] cmd_xbar_demux_003_src3_channel;                                                                        // cmd_xbar_demux_003:src3_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_003_src3_ready;                                                                          // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux_003:src3_ready
	wire          cmd_xbar_demux_003_src5_endofpacket;                                                                    // cmd_xbar_demux_003:src5_endofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_003_src5_valid;                                                                          // cmd_xbar_demux_003:src5_valid -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_003_src5_startofpacket;                                                                  // cmd_xbar_demux_003:src5_startofpacket -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src5_data;                                                                           // cmd_xbar_demux_003:src5_data -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_demux_003_src5_channel;                                                                        // cmd_xbar_demux_003:src5_channel -> dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                    // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_001:sink2_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                          // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_001:sink2_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                                  // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_001:sink2_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src0_data;                                                                           // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_001:sink2_data
	wire    [5:0] cmd_xbar_demux_004_src0_channel;                                                                        // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_001:sink2_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                          // cmd_xbar_mux_001:sink2_ready -> cmd_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_004_src2_endofpacket;                                                                    // cmd_xbar_demux_004:src2_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_004_src2_valid;                                                                          // cmd_xbar_demux_004:src2_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_004_src2_startofpacket;                                                                  // cmd_xbar_demux_004:src2_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src2_data;                                                                           // cmd_xbar_demux_004:src2_data -> cmd_xbar_mux_004:sink1_data
	wire    [5:0] cmd_xbar_demux_004_src2_channel;                                                                        // cmd_xbar_demux_004:src2_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_004_src2_ready;                                                                          // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_004:src2_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                    // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_003:sink2_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                          // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_003:sink2_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                                  // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_003:sink2_startofpacket
	wire  [214:0] cmd_xbar_demux_005_src0_data;                                                                           // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_003:sink2_data
	wire    [5:0] cmd_xbar_demux_005_src0_channel;                                                                        // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_003:sink2_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                          // cmd_xbar_mux_003:sink2_ready -> cmd_xbar_demux_005:src0_ready
	wire          cmd_xbar_demux_006_src0_endofpacket;                                                                    // cmd_xbar_demux_006:src0_endofpacket -> cmd_xbar_mux_005:sink2_endofpacket
	wire          cmd_xbar_demux_006_src0_valid;                                                                          // cmd_xbar_demux_006:src0_valid -> cmd_xbar_mux_005:sink2_valid
	wire          cmd_xbar_demux_006_src0_startofpacket;                                                                  // cmd_xbar_demux_006:src0_startofpacket -> cmd_xbar_mux_005:sink2_startofpacket
	wire  [214:0] cmd_xbar_demux_006_src0_data;                                                                           // cmd_xbar_demux_006:src0_data -> cmd_xbar_mux_005:sink2_data
	wire    [5:0] cmd_xbar_demux_006_src0_channel;                                                                        // cmd_xbar_demux_006:src0_channel -> cmd_xbar_mux_005:sink2_channel
	wire          cmd_xbar_demux_006_src0_ready;                                                                          // cmd_xbar_mux_005:sink2_ready -> cmd_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_001_src1_endofpacket;                                                                    // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_003:sink0_endofpacket
	wire          rsp_xbar_demux_001_src1_valid;                                                                          // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_003:sink0_valid
	wire          rsp_xbar_demux_001_src1_startofpacket;                                                                  // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_003:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src1_data;                                                                           // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_003:sink0_data
	wire    [5:0] rsp_xbar_demux_001_src1_channel;                                                                        // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_003:sink0_channel
	wire          rsp_xbar_demux_001_src1_ready;                                                                          // rsp_xbar_mux_003:sink0_ready -> rsp_xbar_demux_001:src1_ready
	wire          rsp_xbar_demux_001_src2_endofpacket;                                                                    // rsp_xbar_demux_001:src2_endofpacket -> rsp_xbar_mux_004:sink0_endofpacket
	wire          rsp_xbar_demux_001_src2_valid;                                                                          // rsp_xbar_demux_001:src2_valid -> rsp_xbar_mux_004:sink0_valid
	wire          rsp_xbar_demux_001_src2_startofpacket;                                                                  // rsp_xbar_demux_001:src2_startofpacket -> rsp_xbar_mux_004:sink0_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src2_data;                                                                           // rsp_xbar_demux_001:src2_data -> rsp_xbar_mux_004:sink0_data
	wire    [5:0] rsp_xbar_demux_001_src2_channel;                                                                        // rsp_xbar_demux_001:src2_channel -> rsp_xbar_mux_004:sink0_channel
	wire          rsp_xbar_demux_001_src2_ready;                                                                          // rsp_xbar_mux_004:sink0_ready -> rsp_xbar_demux_001:src2_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                    // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_003:sink1_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                          // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_003:sink1_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                                  // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_003:sink1_startofpacket
	wire  [106:0] rsp_xbar_demux_002_src0_data;                                                                           // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_003:sink1_data
	wire    [5:0] rsp_xbar_demux_002_src0_channel;                                                                        // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_003:sink1_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                          // rsp_xbar_mux_003:sink1_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src2_endofpacket;                                                                    // rsp_xbar_demux_003:src2_endofpacket -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_003_src2_valid;                                                                          // rsp_xbar_demux_003:src2_valid -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_003_src2_startofpacket;                                                                  // rsp_xbar_demux_003:src2_startofpacket -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [214:0] rsp_xbar_demux_003_src2_data;                                                                           // rsp_xbar_demux_003:src2_data -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] rsp_xbar_demux_003_src2_channel;                                                                        // rsp_xbar_demux_003:src2_channel -> dma_0_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                    // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_003:sink3_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                          // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_003:sink3_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                                  // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_003:sink3_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src0_data;                                                                           // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_003:sink3_data
	wire    [5:0] rsp_xbar_demux_004_src0_channel;                                                                        // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_003:sink3_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                          // rsp_xbar_mux_003:sink3_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                    // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_004:sink2_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                          // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_004:sink2_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                                  // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_004:sink2_startofpacket
	wire  [106:0] rsp_xbar_demux_004_src1_data;                                                                           // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_004:sink2_data
	wire    [5:0] rsp_xbar_demux_004_src1_channel;                                                                        // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_004:sink2_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                          // rsp_xbar_mux_004:sink2_ready -> rsp_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_005_src2_endofpacket;                                                                    // rsp_xbar_demux_005:src2_endofpacket -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_005_src2_valid;                                                                          // rsp_xbar_demux_005:src2_valid -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_005_src2_startofpacket;                                                                  // rsp_xbar_demux_005:src2_startofpacket -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [214:0] rsp_xbar_demux_005_src2_data;                                                                           // rsp_xbar_demux_005:src2_data -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] rsp_xbar_demux_005_src2_channel;                                                                        // rsp_xbar_demux_005:src2_channel -> dma_0_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                    // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_003:sink5_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                          // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_003:sink5_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                                  // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_003:sink5_startofpacket
	wire  [106:0] rsp_xbar_demux_006_src0_data;                                                                           // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_003:sink5_data
	wire    [5:0] rsp_xbar_demux_006_src0_channel;                                                                        // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_003:sink5_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                          // rsp_xbar_mux_003:sink5_ready -> rsp_xbar_demux_006:src0_ready
	wire          addr_router_002_src_endofpacket;                                                                        // addr_router_002:src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          addr_router_002_src_valid;                                                                              // addr_router_002:src_valid -> cmd_xbar_demux_002:sink_valid
	wire          addr_router_002_src_startofpacket;                                                                      // addr_router_002:src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [106:0] addr_router_002_src_data;                                                                               // addr_router_002:src_data -> cmd_xbar_demux_002:sink_data
	wire    [5:0] addr_router_002_src_channel;                                                                            // addr_router_002:src_channel -> cmd_xbar_demux_002:sink_channel
	wire          addr_router_002_src_ready;                                                                              // cmd_xbar_demux_002:sink_ready -> addr_router_002:src_ready
	wire          crosser_003_out_ready;                                                                                  // fir_dma_read_master_translator_avalon_universal_master_0_agent:rp_ready -> crosser_003:out_ready
	wire          limiter_cmd_src_endofpacket;                                                                            // limiter:cmd_src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                          // limiter:cmd_src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [106:0] limiter_cmd_src_data;                                                                                   // limiter:cmd_src_data -> cmd_xbar_demux_003:sink_data
	wire    [5:0] limiter_cmd_src_channel;                                                                                // limiter:cmd_src_channel -> cmd_xbar_demux_003:sink_channel
	wire          limiter_cmd_src_ready;                                                                                  // cmd_xbar_demux_003:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_003_src_endofpacket;                                                                       // rsp_xbar_mux_003:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_003_src_valid;                                                                             // rsp_xbar_mux_003:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_003_src_startofpacket;                                                                     // rsp_xbar_mux_003:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_003_src_data;                                                                              // rsp_xbar_mux_003:src_data -> limiter:rsp_sink_data
	wire    [5:0] rsp_xbar_mux_003_src_channel;                                                                           // rsp_xbar_mux_003:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_003_src_ready;                                                                             // limiter:rsp_sink_ready -> rsp_xbar_mux_003:src_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                        // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                      // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [106:0] limiter_001_cmd_src_data;                                                                               // limiter_001:cmd_src_data -> cmd_xbar_demux_004:sink_data
	wire    [5:0] limiter_001_cmd_src_channel;                                                                            // limiter_001:cmd_src_channel -> cmd_xbar_demux_004:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                              // cmd_xbar_demux_004:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_004_src_endofpacket;                                                                       // rsp_xbar_mux_004:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_004_src_valid;                                                                             // rsp_xbar_mux_004:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_004_src_startofpacket;                                                                     // rsp_xbar_mux_004:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [106:0] rsp_xbar_mux_004_src_data;                                                                              // rsp_xbar_mux_004:src_data -> limiter_001:rsp_sink_data
	wire    [5:0] rsp_xbar_mux_004_src_channel;                                                                           // rsp_xbar_mux_004:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_004_src_ready;                                                                             // limiter_001:rsp_sink_ready -> rsp_xbar_mux_004:src_ready
	wire          addr_router_005_src_endofpacket;                                                                        // addr_router_005:src_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          addr_router_005_src_valid;                                                                              // addr_router_005:src_valid -> cmd_xbar_demux_005:sink_valid
	wire          addr_router_005_src_startofpacket;                                                                      // addr_router_005:src_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [214:0] addr_router_005_src_data;                                                                               // addr_router_005:src_data -> cmd_xbar_demux_005:sink_data
	wire    [5:0] addr_router_005_src_channel;                                                                            // addr_router_005:src_channel -> cmd_xbar_demux_005:sink_channel
	wire          addr_router_005_src_ready;                                                                              // cmd_xbar_demux_005:sink_ready -> addr_router_005:src_ready
	wire          rsp_xbar_demux_003_src2_ready;                                                                          // dma_0_read_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_003:src2_ready
	wire          addr_router_006_src_endofpacket;                                                                        // addr_router_006:src_endofpacket -> cmd_xbar_demux_006:sink_endofpacket
	wire          addr_router_006_src_valid;                                                                              // addr_router_006:src_valid -> cmd_xbar_demux_006:sink_valid
	wire          addr_router_006_src_startofpacket;                                                                      // addr_router_006:src_startofpacket -> cmd_xbar_demux_006:sink_startofpacket
	wire  [214:0] addr_router_006_src_data;                                                                               // addr_router_006:src_data -> cmd_xbar_demux_006:sink_data
	wire    [5:0] addr_router_006_src_channel;                                                                            // addr_router_006:src_channel -> cmd_xbar_demux_006:sink_channel
	wire          addr_router_006_src_ready;                                                                              // cmd_xbar_demux_006:sink_ready -> addr_router_006:src_ready
	wire          rsp_xbar_demux_005_src2_ready;                                                                          // dma_0_write_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_005:src2_ready
	wire          cmd_xbar_mux_001_src_endofpacket;                                                                       // cmd_xbar_mux_001:src_endofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_001_src_valid;                                                                             // cmd_xbar_mux_001:src_valid -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_001_src_startofpacket;                                                                     // cmd_xbar_mux_001:src_startofpacket -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_001_src_data;                                                                              // cmd_xbar_mux_001:src_data -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_001_src_channel;                                                                           // cmd_xbar_mux_001:src_channel -> flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_001_src_ready;                                                                             // flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire          id_router_001_src_endofpacket;                                                                          // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          id_router_001_src_valid;                                                                                // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire          id_router_001_src_startofpacket;                                                                        // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [106:0] id_router_001_src_data;                                                                                 // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire    [5:0] id_router_001_src_channel;                                                                              // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire          id_router_001_src_ready;                                                                                // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire          cmd_xbar_demux_003_src1_ready;                                                                          // slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src1_ready
	wire          id_router_002_src_endofpacket;                                                                          // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                                // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                        // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [106:0] id_router_002_src_data;                                                                                 // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [5:0] id_router_002_src_channel;                                                                              // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                                // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                       // cmd_xbar_mux_003:src_endofpacket -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                             // cmd_xbar_mux_003:src_valid -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                     // cmd_xbar_mux_003:src_startofpacket -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [214:0] cmd_xbar_mux_003_src_data;                                                                              // cmd_xbar_mux_003:src_data -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_003_src_channel;                                                                           // cmd_xbar_mux_003:src_channel -> ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                             // ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                          // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                                // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                        // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [214:0] id_router_003_src_data;                                                                                 // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [5:0] id_router_003_src_channel;                                                                              // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                                // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                       // cmd_xbar_mux_004:src_endofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                             // cmd_xbar_mux_004:src_valid -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                     // cmd_xbar_mux_004:src_startofpacket -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [106:0] cmd_xbar_mux_004_src_data;                                                                              // cmd_xbar_mux_004:src_data -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_004_src_channel;                                                                           // cmd_xbar_mux_004:src_channel -> cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                             // cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	wire          id_router_004_src_endofpacket;                                                                          // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                                // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                        // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [106:0] id_router_004_src_data;                                                                                 // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [5:0] id_router_004_src_channel;                                                                              // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                                // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                       // cmd_xbar_mux_005:src_endofpacket -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                             // cmd_xbar_mux_005:src_valid -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                     // cmd_xbar_mux_005:src_startofpacket -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [214:0] cmd_xbar_mux_005_src_data;                                                                              // cmd_xbar_mux_005:src_data -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_data
	wire    [5:0] cmd_xbar_mux_005_src_channel;                                                                           // cmd_xbar_mux_005:src_channel -> ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                             // ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                          // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                                // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                        // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [214:0] id_router_005_src_data;                                                                                 // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [5:0] id_router_005_src_channel;                                                                              // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                                // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_demux_003_src5_ready;                                                                          // dma_0_control_port_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_003:src5_ready
	wire          id_router_006_src_endofpacket;                                                                          // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                                // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                        // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [106:0] id_router_006_src_data;                                                                                 // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [5:0] id_router_006_src_channel;                                                                              // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                                // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_demux_007_src0_endofpacket;                                                                    // cmd_xbar_demux_007:src0_endofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src0_valid;                                                                          // cmd_xbar_demux_007:src0_valid -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src0_startofpacket;                                                                  // cmd_xbar_demux_007:src0_startofpacket -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src0_data;                                                                           // cmd_xbar_demux_007:src0_data -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src0_channel;                                                                        // cmd_xbar_demux_007:src0_channel -> high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src1_endofpacket;                                                                    // cmd_xbar_demux_007:src1_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src1_valid;                                                                          // cmd_xbar_demux_007:src1_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src1_startofpacket;                                                                  // cmd_xbar_demux_007:src1_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src1_data;                                                                           // cmd_xbar_demux_007:src1_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src1_channel;                                                                        // cmd_xbar_demux_007:src1_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src2_endofpacket;                                                                    // cmd_xbar_demux_007:src2_endofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src2_valid;                                                                          // cmd_xbar_demux_007:src2_valid -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src2_startofpacket;                                                                  // cmd_xbar_demux_007:src2_startofpacket -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src2_data;                                                                           // cmd_xbar_demux_007:src2_data -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src2_channel;                                                                        // cmd_xbar_demux_007:src2_channel -> performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src3_endofpacket;                                                                    // cmd_xbar_demux_007:src3_endofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src3_valid;                                                                          // cmd_xbar_demux_007:src3_valid -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src3_startofpacket;                                                                  // cmd_xbar_demux_007:src3_startofpacket -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src3_data;                                                                           // cmd_xbar_demux_007:src3_data -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src3_channel;                                                                        // cmd_xbar_demux_007:src3_channel -> sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src4_endofpacket;                                                                    // cmd_xbar_demux_007:src4_endofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src4_valid;                                                                          // cmd_xbar_demux_007:src4_valid -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src4_startofpacket;                                                                  // cmd_xbar_demux_007:src4_startofpacket -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src4_data;                                                                           // cmd_xbar_demux_007:src4_data -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src4_channel;                                                                        // cmd_xbar_demux_007:src4_channel -> sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src7_endofpacket;                                                                    // cmd_xbar_demux_007:src7_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src7_valid;                                                                          // cmd_xbar_demux_007:src7_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src7_startofpacket;                                                                  // cmd_xbar_demux_007:src7_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src7_data;                                                                           // cmd_xbar_demux_007:src7_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src7_channel;                                                                        // cmd_xbar_demux_007:src7_channel -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src8_endofpacket;                                                                    // cmd_xbar_demux_007:src8_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src8_valid;                                                                          // cmd_xbar_demux_007:src8_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src8_startofpacket;                                                                  // cmd_xbar_demux_007:src8_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src8_data;                                                                           // cmd_xbar_demux_007:src8_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src8_channel;                                                                        // cmd_xbar_demux_007:src8_channel -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src9_endofpacket;                                                                    // cmd_xbar_demux_007:src9_endofpacket -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src9_valid;                                                                          // cmd_xbar_demux_007:src9_valid -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src9_startofpacket;                                                                  // cmd_xbar_demux_007:src9_startofpacket -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src9_data;                                                                           // cmd_xbar_demux_007:src9_data -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src9_channel;                                                                        // cmd_xbar_demux_007:src9_channel -> lcd_display_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src10_endofpacket;                                                                   // cmd_xbar_demux_007:src10_endofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_007_src10_valid;                                                                         // cmd_xbar_demux_007:src10_valid -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_007_src10_startofpacket;                                                                 // cmd_xbar_demux_007:src10_startofpacket -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src10_data;                                                                          // cmd_xbar_demux_007:src10_data -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] cmd_xbar_demux_007_src10_channel;                                                                       // cmd_xbar_demux_007:src10_channel -> seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                    // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_007:sink0_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                          // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_007:sink0_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                                  // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_007:sink0_startofpacket
	wire   [82:0] rsp_xbar_demux_007_src0_data;                                                                           // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_007:sink0_data
	wire   [10:0] rsp_xbar_demux_007_src0_channel;                                                                        // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_007:sink0_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                          // rsp_xbar_mux_007:sink0_ready -> rsp_xbar_demux_007:src0_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                    // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_007:sink1_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                          // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_007:sink1_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                                  // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_007:sink1_startofpacket
	wire   [82:0] rsp_xbar_demux_008_src0_data;                                                                           // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_007:sink1_data
	wire   [10:0] rsp_xbar_demux_008_src0_channel;                                                                        // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_007:sink1_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                          // rsp_xbar_mux_007:sink1_ready -> rsp_xbar_demux_008:src0_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                    // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_007:sink2_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                          // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_007:sink2_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                                  // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_007:sink2_startofpacket
	wire   [82:0] rsp_xbar_demux_009_src0_data;                                                                           // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_007:sink2_data
	wire   [10:0] rsp_xbar_demux_009_src0_channel;                                                                        // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_007:sink2_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                          // rsp_xbar_mux_007:sink2_ready -> rsp_xbar_demux_009:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                    // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_007:sink3_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                          // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_007:sink3_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                                  // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_007:sink3_startofpacket
	wire   [82:0] rsp_xbar_demux_010_src0_data;                                                                           // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_007:sink3_data
	wire   [10:0] rsp_xbar_demux_010_src0_channel;                                                                        // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_007:sink3_channel
	wire          rsp_xbar_demux_010_src0_ready;                                                                          // rsp_xbar_mux_007:sink3_ready -> rsp_xbar_demux_010:src0_ready
	wire          rsp_xbar_demux_011_src0_endofpacket;                                                                    // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_007:sink4_endofpacket
	wire          rsp_xbar_demux_011_src0_valid;                                                                          // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_007:sink4_valid
	wire          rsp_xbar_demux_011_src0_startofpacket;                                                                  // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_007:sink4_startofpacket
	wire   [82:0] rsp_xbar_demux_011_src0_data;                                                                           // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_007:sink4_data
	wire   [10:0] rsp_xbar_demux_011_src0_channel;                                                                        // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_007:sink4_channel
	wire          rsp_xbar_demux_011_src0_ready;                                                                          // rsp_xbar_mux_007:sink4_ready -> rsp_xbar_demux_011:src0_ready
	wire          rsp_xbar_demux_014_src0_endofpacket;                                                                    // rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_007:sink7_endofpacket
	wire          rsp_xbar_demux_014_src0_valid;                                                                          // rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_007:sink7_valid
	wire          rsp_xbar_demux_014_src0_startofpacket;                                                                  // rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_007:sink7_startofpacket
	wire   [82:0] rsp_xbar_demux_014_src0_data;                                                                           // rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_007:sink7_data
	wire   [10:0] rsp_xbar_demux_014_src0_channel;                                                                        // rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_007:sink7_channel
	wire          rsp_xbar_demux_014_src0_ready;                                                                          // rsp_xbar_mux_007:sink7_ready -> rsp_xbar_demux_014:src0_ready
	wire          rsp_xbar_demux_015_src0_endofpacket;                                                                    // rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_007:sink8_endofpacket
	wire          rsp_xbar_demux_015_src0_valid;                                                                          // rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_007:sink8_valid
	wire          rsp_xbar_demux_015_src0_startofpacket;                                                                  // rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_007:sink8_startofpacket
	wire   [82:0] rsp_xbar_demux_015_src0_data;                                                                           // rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_007:sink8_data
	wire   [10:0] rsp_xbar_demux_015_src0_channel;                                                                        // rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_007:sink8_channel
	wire          rsp_xbar_demux_015_src0_ready;                                                                          // rsp_xbar_mux_007:sink8_ready -> rsp_xbar_demux_015:src0_ready
	wire          rsp_xbar_demux_016_src0_endofpacket;                                                                    // rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_007:sink9_endofpacket
	wire          rsp_xbar_demux_016_src0_valid;                                                                          // rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_007:sink9_valid
	wire          rsp_xbar_demux_016_src0_startofpacket;                                                                  // rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_007:sink9_startofpacket
	wire   [82:0] rsp_xbar_demux_016_src0_data;                                                                           // rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_007:sink9_data
	wire   [10:0] rsp_xbar_demux_016_src0_channel;                                                                        // rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_007:sink9_channel
	wire          rsp_xbar_demux_016_src0_ready;                                                                          // rsp_xbar_mux_007:sink9_ready -> rsp_xbar_demux_016:src0_ready
	wire          rsp_xbar_demux_017_src0_endofpacket;                                                                    // rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_007:sink10_endofpacket
	wire          rsp_xbar_demux_017_src0_valid;                                                                          // rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_007:sink10_valid
	wire          rsp_xbar_demux_017_src0_startofpacket;                                                                  // rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_007:sink10_startofpacket
	wire   [82:0] rsp_xbar_demux_017_src0_data;                                                                           // rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_007:sink10_data
	wire   [10:0] rsp_xbar_demux_017_src0_channel;                                                                        // rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_007:sink10_channel
	wire          rsp_xbar_demux_017_src0_ready;                                                                          // rsp_xbar_mux_007:sink10_ready -> rsp_xbar_demux_017:src0_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                        // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_007:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                      // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_007:sink_startofpacket
	wire   [82:0] limiter_002_cmd_src_data;                                                                               // limiter_002:cmd_src_data -> cmd_xbar_demux_007:sink_data
	wire   [10:0] limiter_002_cmd_src_channel;                                                                            // limiter_002:cmd_src_channel -> cmd_xbar_demux_007:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                              // cmd_xbar_demux_007:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_007_src_endofpacket;                                                                       // rsp_xbar_mux_007:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_007_src_valid;                                                                             // rsp_xbar_mux_007:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_007_src_startofpacket;                                                                     // rsp_xbar_mux_007:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire   [82:0] rsp_xbar_mux_007_src_data;                                                                              // rsp_xbar_mux_007:src_data -> limiter_002:rsp_sink_data
	wire   [10:0] rsp_xbar_mux_007_src_channel;                                                                           // rsp_xbar_mux_007:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_007_src_ready;                                                                             // limiter_002:rsp_sink_ready -> rsp_xbar_mux_007:src_ready
	wire          cmd_xbar_demux_007_src0_ready;                                                                          // high_res_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src0_ready
	wire          id_router_007_src_endofpacket;                                                                          // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                                // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                        // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire   [82:0] id_router_007_src_data;                                                                                 // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire   [10:0] id_router_007_src_channel;                                                                              // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                                // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_demux_007_src1_ready;                                                                          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src1_ready
	wire          id_router_008_src_endofpacket;                                                                          // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                                // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                        // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire   [82:0] id_router_008_src_data;                                                                                 // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire   [10:0] id_router_008_src_channel;                                                                              // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                                // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_demux_007_src2_ready;                                                                          // performance_counter_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src2_ready
	wire          id_router_009_src_endofpacket;                                                                          // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                                // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                        // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire   [82:0] id_router_009_src_data;                                                                                 // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire   [10:0] id_router_009_src_channel;                                                                              // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                                // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_007_src3_ready;                                                                          // sys_clk_timer_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src3_ready
	wire          id_router_010_src_endofpacket;                                                                          // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          id_router_010_src_valid;                                                                                // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire          id_router_010_src_startofpacket;                                                                        // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire   [82:0] id_router_010_src_data;                                                                                 // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire   [10:0] id_router_010_src_channel;                                                                              // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire          id_router_010_src_ready;                                                                                // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire          cmd_xbar_demux_007_src4_ready;                                                                          // sysid_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src4_ready
	wire          id_router_011_src_endofpacket;                                                                          // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire          id_router_011_src_valid;                                                                                // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire          id_router_011_src_startofpacket;                                                                        // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire   [82:0] id_router_011_src_data;                                                                                 // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire   [10:0] id_router_011_src_channel;                                                                              // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire          id_router_011_src_ready;                                                                                // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire          crosser_004_out_ready;                                                                                  // fir_dma_control_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_004:out_ready
	wire          id_router_012_src_endofpacket;                                                                          // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire          id_router_012_src_valid;                                                                                // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire          id_router_012_src_startofpacket;                                                                        // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire   [82:0] id_router_012_src_data;                                                                                 // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire   [10:0] id_router_012_src_channel;                                                                              // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire          id_router_012_src_ready;                                                                                // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire          crosser_005_out_ready;                                                                                  // pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_ready -> crosser_005:out_ready
	wire          id_router_013_src_endofpacket;                                                                          // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire          id_router_013_src_valid;                                                                                // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire          id_router_013_src_startofpacket;                                                                        // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire   [82:0] id_router_013_src_data;                                                                                 // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire   [10:0] id_router_013_src_channel;                                                                              // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire          id_router_013_src_ready;                                                                                // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire          cmd_xbar_demux_007_src7_ready;                                                                          // button_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src7_ready
	wire          id_router_014_src_endofpacket;                                                                          // id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	wire          id_router_014_src_valid;                                                                                // id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	wire          id_router_014_src_startofpacket;                                                                        // id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	wire   [82:0] id_router_014_src_data;                                                                                 // id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	wire   [10:0] id_router_014_src_channel;                                                                              // id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	wire          id_router_014_src_ready;                                                                                // rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	wire          cmd_xbar_demux_007_src8_ready;                                                                          // led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src8_ready
	wire          id_router_015_src_endofpacket;                                                                          // id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	wire          id_router_015_src_valid;                                                                                // id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	wire          id_router_015_src_startofpacket;                                                                        // id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	wire   [82:0] id_router_015_src_data;                                                                                 // id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	wire   [10:0] id_router_015_src_channel;                                                                              // id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	wire          id_router_015_src_ready;                                                                                // rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	wire          cmd_xbar_demux_007_src9_ready;                                                                          // lcd_display_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src9_ready
	wire          id_router_016_src_endofpacket;                                                                          // id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	wire          id_router_016_src_valid;                                                                                // id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	wire          id_router_016_src_startofpacket;                                                                        // id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	wire   [82:0] id_router_016_src_data;                                                                                 // id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	wire   [10:0] id_router_016_src_channel;                                                                              // id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	wire          id_router_016_src_ready;                                                                                // rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	wire          cmd_xbar_demux_007_src10_ready;                                                                         // seven_seg_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_007:src10_ready
	wire          id_router_017_src_endofpacket;                                                                          // id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	wire          id_router_017_src_valid;                                                                                // id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	wire          id_router_017_src_startofpacket;                                                                        // id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	wire   [82:0] id_router_017_src_data;                                                                                 // id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	wire   [10:0] id_router_017_src_channel;                                                                              // id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	wire          id_router_017_src_ready;                                                                                // rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	wire          cmd_xbar_demux_008_src0_endofpacket;                                                                    // cmd_xbar_demux_008:src0_endofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_008_src0_valid;                                                                          // cmd_xbar_demux_008:src0_valid -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_008_src0_startofpacket;                                                                  // cmd_xbar_demux_008:src0_startofpacket -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [93:0] cmd_xbar_demux_008_src0_data;                                                                           // cmd_xbar_demux_008:src0_data -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_data
	wire    [1:0] cmd_xbar_demux_008_src0_channel;                                                                        // cmd_xbar_demux_008:src0_channel -> ssram_uas_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_008_src1_endofpacket;                                                                    // cmd_xbar_demux_008:src1_endofpacket -> width_adapter_012:in_endofpacket
	wire          cmd_xbar_demux_008_src1_valid;                                                                          // cmd_xbar_demux_008:src1_valid -> width_adapter_012:in_valid
	wire          cmd_xbar_demux_008_src1_startofpacket;                                                                  // cmd_xbar_demux_008:src1_startofpacket -> width_adapter_012:in_startofpacket
	wire   [93:0] cmd_xbar_demux_008_src1_data;                                                                           // cmd_xbar_demux_008:src1_data -> width_adapter_012:in_data
	wire    [1:0] cmd_xbar_demux_008_src1_channel;                                                                        // cmd_xbar_demux_008:src1_channel -> width_adapter_012:in_channel
	wire          rsp_xbar_demux_018_src0_endofpacket;                                                                    // rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_008:sink0_endofpacket
	wire          rsp_xbar_demux_018_src0_valid;                                                                          // rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_008:sink0_valid
	wire          rsp_xbar_demux_018_src0_startofpacket;                                                                  // rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_008:sink0_startofpacket
	wire   [93:0] rsp_xbar_demux_018_src0_data;                                                                           // rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_008:sink0_data
	wire    [1:0] rsp_xbar_demux_018_src0_channel;                                                                        // rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_008:sink0_channel
	wire          rsp_xbar_demux_018_src0_ready;                                                                          // rsp_xbar_mux_008:sink0_ready -> rsp_xbar_demux_018:src0_ready
	wire          rsp_xbar_demux_019_src0_endofpacket;                                                                    // rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_008:sink1_endofpacket
	wire          rsp_xbar_demux_019_src0_valid;                                                                          // rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_008:sink1_valid
	wire          rsp_xbar_demux_019_src0_startofpacket;                                                                  // rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_008:sink1_startofpacket
	wire   [93:0] rsp_xbar_demux_019_src0_data;                                                                           // rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_008:sink1_data
	wire    [1:0] rsp_xbar_demux_019_src0_channel;                                                                        // rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_008:sink1_channel
	wire          rsp_xbar_demux_019_src0_ready;                                                                          // rsp_xbar_mux_008:sink1_ready -> rsp_xbar_demux_019:src0_ready
	wire          limiter_003_cmd_src_endofpacket;                                                                        // limiter_003:cmd_src_endofpacket -> cmd_xbar_demux_008:sink_endofpacket
	wire          limiter_003_cmd_src_startofpacket;                                                                      // limiter_003:cmd_src_startofpacket -> cmd_xbar_demux_008:sink_startofpacket
	wire   [93:0] limiter_003_cmd_src_data;                                                                               // limiter_003:cmd_src_data -> cmd_xbar_demux_008:sink_data
	wire    [1:0] limiter_003_cmd_src_channel;                                                                            // limiter_003:cmd_src_channel -> cmd_xbar_demux_008:sink_channel
	wire          limiter_003_cmd_src_ready;                                                                              // cmd_xbar_demux_008:sink_ready -> limiter_003:cmd_src_ready
	wire          rsp_xbar_mux_008_src_endofpacket;                                                                       // rsp_xbar_mux_008:src_endofpacket -> limiter_003:rsp_sink_endofpacket
	wire          rsp_xbar_mux_008_src_valid;                                                                             // rsp_xbar_mux_008:src_valid -> limiter_003:rsp_sink_valid
	wire          rsp_xbar_mux_008_src_startofpacket;                                                                     // rsp_xbar_mux_008:src_startofpacket -> limiter_003:rsp_sink_startofpacket
	wire   [93:0] rsp_xbar_mux_008_src_data;                                                                              // rsp_xbar_mux_008:src_data -> limiter_003:rsp_sink_data
	wire    [1:0] rsp_xbar_mux_008_src_channel;                                                                           // rsp_xbar_mux_008:src_channel -> limiter_003:rsp_sink_channel
	wire          rsp_xbar_mux_008_src_ready;                                                                             // limiter_003:rsp_sink_ready -> rsp_xbar_mux_008:src_ready
	wire          cmd_xbar_demux_008_src0_ready;                                                                          // ssram_uas_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_008:src0_ready
	wire          id_router_018_src_endofpacket;                                                                          // id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	wire          id_router_018_src_valid;                                                                                // id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	wire          id_router_018_src_startofpacket;                                                                        // id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	wire   [93:0] id_router_018_src_data;                                                                                 // id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	wire    [1:0] id_router_018_src_channel;                                                                              // id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	wire          id_router_018_src_ready;                                                                                // rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	wire          cmd_xbar_demux_009_src0_endofpacket;                                                                    // cmd_xbar_demux_009:src0_endofpacket -> width_adapter_014:in_endofpacket
	wire          cmd_xbar_demux_009_src0_valid;                                                                          // cmd_xbar_demux_009:src0_valid -> width_adapter_014:in_valid
	wire          cmd_xbar_demux_009_src0_startofpacket;                                                                  // cmd_xbar_demux_009:src0_startofpacket -> width_adapter_014:in_startofpacket
	wire  [204:0] cmd_xbar_demux_009_src0_data;                                                                           // cmd_xbar_demux_009:src0_data -> width_adapter_014:in_data
	wire    [0:0] cmd_xbar_demux_009_src0_channel;                                                                        // cmd_xbar_demux_009:src0_channel -> width_adapter_014:in_channel
	wire          rsp_xbar_demux_020_src0_endofpacket;                                                                    // rsp_xbar_demux_020:src0_endofpacket -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          rsp_xbar_demux_020_src0_valid;                                                                          // rsp_xbar_demux_020:src0_valid -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          rsp_xbar_demux_020_src0_startofpacket;                                                                  // rsp_xbar_demux_020:src0_startofpacket -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [204:0] rsp_xbar_demux_020_src0_data;                                                                           // rsp_xbar_demux_020:src0_data -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire    [0:0] rsp_xbar_demux_020_src0_channel;                                                                        // rsp_xbar_demux_020:src0_channel -> ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_009_src_endofpacket;                                                                        // addr_router_009:src_endofpacket -> cmd_xbar_demux_009:sink_endofpacket
	wire          addr_router_009_src_valid;                                                                              // addr_router_009:src_valid -> cmd_xbar_demux_009:sink_valid
	wire          addr_router_009_src_startofpacket;                                                                      // addr_router_009:src_startofpacket -> cmd_xbar_demux_009:sink_startofpacket
	wire  [204:0] addr_router_009_src_data;                                                                               // addr_router_009:src_data -> cmd_xbar_demux_009:sink_data
	wire    [0:0] addr_router_009_src_channel;                                                                            // addr_router_009:src_channel -> cmd_xbar_demux_009:sink_channel
	wire          addr_router_009_src_ready;                                                                              // cmd_xbar_demux_009:sink_ready -> addr_router_009:src_ready
	wire          rsp_xbar_demux_020_src0_ready;                                                                          // ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_demux_020:src0_ready
	wire          addr_router_src_endofpacket;                                                                            // addr_router:src_endofpacket -> width_adapter:in_endofpacket
	wire          addr_router_src_valid;                                                                                  // addr_router:src_valid -> width_adapter:in_valid
	wire          addr_router_src_startofpacket;                                                                          // addr_router:src_startofpacket -> width_adapter:in_startofpacket
	wire  [101:0] addr_router_src_data;                                                                                   // addr_router:src_data -> width_adapter:in_data
	wire    [1:0] addr_router_src_channel;                                                                                // addr_router:src_channel -> width_adapter:in_channel
	wire          addr_router_src_ready;                                                                                  // width_adapter:in_ready -> addr_router:src_ready
	wire          width_adapter_src_endofpacket;                                                                          // width_adapter:out_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          width_adapter_src_valid;                                                                                // width_adapter:out_valid -> cmd_xbar_demux:sink_valid
	wire          width_adapter_src_startofpacket;                                                                        // width_adapter:out_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [137:0] width_adapter_src_data;                                                                                 // width_adapter:out_data -> cmd_xbar_demux:sink_data
	wire          width_adapter_src_ready;                                                                                // cmd_xbar_demux:sink_ready -> width_adapter:out_ready
	wire    [1:0] width_adapter_src_channel;                                                                              // width_adapter:out_channel -> cmd_xbar_demux:sink_channel
	wire          crosser_001_out_ready;                                                                                  // width_adapter_001:in_ready -> crosser_001:out_ready
	wire          width_adapter_001_src_endofpacket;                                                                      // width_adapter_001:out_endofpacket -> fir_dma_write_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          width_adapter_001_src_valid;                                                                            // width_adapter_001:out_valid -> fir_dma_write_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          width_adapter_001_src_startofpacket;                                                                    // width_adapter_001:out_startofpacket -> fir_dma_write_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [101:0] width_adapter_001_src_data;                                                                             // width_adapter_001:out_data -> fir_dma_write_master_translator_avalon_universal_master_0_agent:rp_data
	wire          width_adapter_001_src_ready;                                                                            // fir_dma_write_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_001:out_ready
	wire    [1:0] width_adapter_001_src_channel;                                                                          // width_adapter_001:out_channel -> fir_dma_write_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          addr_router_001_src_endofpacket;                                                                        // addr_router_001:src_endofpacket -> width_adapter_002:in_endofpacket
	wire          addr_router_001_src_valid;                                                                              // addr_router_001:src_valid -> width_adapter_002:in_valid
	wire          addr_router_001_src_startofpacket;                                                                      // addr_router_001:src_startofpacket -> width_adapter_002:in_startofpacket
	wire  [209:0] addr_router_001_src_data;                                                                               // addr_router_001:src_data -> width_adapter_002:in_data
	wire    [1:0] addr_router_001_src_channel;                                                                            // addr_router_001:src_channel -> width_adapter_002:in_channel
	wire          addr_router_001_src_ready;                                                                              // width_adapter_002:in_ready -> addr_router_001:src_ready
	wire          width_adapter_002_src_endofpacket;                                                                      // width_adapter_002:out_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          width_adapter_002_src_valid;                                                                            // width_adapter_002:out_valid -> cmd_xbar_demux_001:sink_valid
	wire          width_adapter_002_src_startofpacket;                                                                    // width_adapter_002:out_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [137:0] width_adapter_002_src_data;                                                                             // width_adapter_002:out_data -> cmd_xbar_demux_001:sink_data
	wire          width_adapter_002_src_ready;                                                                            // cmd_xbar_demux_001:sink_ready -> width_adapter_002:out_ready
	wire    [1:0] width_adapter_002_src_channel;                                                                          // width_adapter_002:out_channel -> cmd_xbar_demux_001:sink_channel
	wire          rsp_xbar_demux_src1_ready;                                                                              // width_adapter_003:in_ready -> rsp_xbar_demux:src1_ready
	wire          width_adapter_003_src_endofpacket;                                                                      // width_adapter_003:out_endofpacket -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          width_adapter_003_src_valid;                                                                            // width_adapter_003:out_valid -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_valid
	wire          width_adapter_003_src_startofpacket;                                                                    // width_adapter_003:out_startofpacket -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [209:0] width_adapter_003_src_data;                                                                             // width_adapter_003:out_data -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_data
	wire          width_adapter_003_src_ready;                                                                            // ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_003:out_ready
	wire    [1:0] width_adapter_003_src_channel;                                                                          // width_adapter_003:out_channel -> ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent:rp_channel
	wire          cmd_xbar_demux_003_src2_endofpacket;                                                                    // cmd_xbar_demux_003:src2_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_003_src2_valid;                                                                          // cmd_xbar_demux_003:src2_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_003_src2_startofpacket;                                                                  // cmd_xbar_demux_003:src2_startofpacket -> width_adapter_004:in_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src2_data;                                                                           // cmd_xbar_demux_003:src2_data -> width_adapter_004:in_data
	wire    [5:0] cmd_xbar_demux_003_src2_channel;                                                                        // cmd_xbar_demux_003:src2_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_003_src2_ready;                                                                          // width_adapter_004:in_ready -> cmd_xbar_demux_003:src2_ready
	wire          width_adapter_004_src_endofpacket;                                                                      // width_adapter_004:out_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                                            // width_adapter_004:out_valid -> cmd_xbar_mux_003:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                                    // width_adapter_004:out_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [214:0] width_adapter_004_src_data;                                                                             // width_adapter_004:out_data -> cmd_xbar_mux_003:sink0_data
	wire          width_adapter_004_src_ready;                                                                            // cmd_xbar_mux_003:sink0_ready -> width_adapter_004:out_ready
	wire    [5:0] width_adapter_004_src_channel;                                                                          // width_adapter_004:out_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_003_src4_endofpacket;                                                                    // cmd_xbar_demux_003:src4_endofpacket -> width_adapter_005:in_endofpacket
	wire          cmd_xbar_demux_003_src4_valid;                                                                          // cmd_xbar_demux_003:src4_valid -> width_adapter_005:in_valid
	wire          cmd_xbar_demux_003_src4_startofpacket;                                                                  // cmd_xbar_demux_003:src4_startofpacket -> width_adapter_005:in_startofpacket
	wire  [106:0] cmd_xbar_demux_003_src4_data;                                                                           // cmd_xbar_demux_003:src4_data -> width_adapter_005:in_data
	wire    [5:0] cmd_xbar_demux_003_src4_channel;                                                                        // cmd_xbar_demux_003:src4_channel -> width_adapter_005:in_channel
	wire          cmd_xbar_demux_003_src4_ready;                                                                          // width_adapter_005:in_ready -> cmd_xbar_demux_003:src4_ready
	wire          width_adapter_005_src_endofpacket;                                                                      // width_adapter_005:out_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          width_adapter_005_src_valid;                                                                            // width_adapter_005:out_valid -> cmd_xbar_mux_005:sink0_valid
	wire          width_adapter_005_src_startofpacket;                                                                    // width_adapter_005:out_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [214:0] width_adapter_005_src_data;                                                                             // width_adapter_005:out_data -> cmd_xbar_mux_005:sink0_data
	wire          width_adapter_005_src_ready;                                                                            // cmd_xbar_mux_005:sink0_ready -> width_adapter_005:out_ready
	wire    [5:0] width_adapter_005_src_channel;                                                                          // width_adapter_005:out_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_004_src1_endofpacket;                                                                    // cmd_xbar_demux_004:src1_endofpacket -> width_adapter_006:in_endofpacket
	wire          cmd_xbar_demux_004_src1_valid;                                                                          // cmd_xbar_demux_004:src1_valid -> width_adapter_006:in_valid
	wire          cmd_xbar_demux_004_src1_startofpacket;                                                                  // cmd_xbar_demux_004:src1_startofpacket -> width_adapter_006:in_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src1_data;                                                                           // cmd_xbar_demux_004:src1_data -> width_adapter_006:in_data
	wire    [5:0] cmd_xbar_demux_004_src1_channel;                                                                        // cmd_xbar_demux_004:src1_channel -> width_adapter_006:in_channel
	wire          cmd_xbar_demux_004_src1_ready;                                                                          // width_adapter_006:in_ready -> cmd_xbar_demux_004:src1_ready
	wire          width_adapter_006_src_endofpacket;                                                                      // width_adapter_006:out_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          width_adapter_006_src_valid;                                                                            // width_adapter_006:out_valid -> cmd_xbar_mux_003:sink1_valid
	wire          width_adapter_006_src_startofpacket;                                                                    // width_adapter_006:out_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [214:0] width_adapter_006_src_data;                                                                             // width_adapter_006:out_data -> cmd_xbar_mux_003:sink1_data
	wire          width_adapter_006_src_ready;                                                                            // cmd_xbar_mux_003:sink1_ready -> width_adapter_006:out_ready
	wire    [5:0] width_adapter_006_src_channel;                                                                          // width_adapter_006:out_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_004_src3_endofpacket;                                                                    // cmd_xbar_demux_004:src3_endofpacket -> width_adapter_007:in_endofpacket
	wire          cmd_xbar_demux_004_src3_valid;                                                                          // cmd_xbar_demux_004:src3_valid -> width_adapter_007:in_valid
	wire          cmd_xbar_demux_004_src3_startofpacket;                                                                  // cmd_xbar_demux_004:src3_startofpacket -> width_adapter_007:in_startofpacket
	wire  [106:0] cmd_xbar_demux_004_src3_data;                                                                           // cmd_xbar_demux_004:src3_data -> width_adapter_007:in_data
	wire    [5:0] cmd_xbar_demux_004_src3_channel;                                                                        // cmd_xbar_demux_004:src3_channel -> width_adapter_007:in_channel
	wire          cmd_xbar_demux_004_src3_ready;                                                                          // width_adapter_007:in_ready -> cmd_xbar_demux_004:src3_ready
	wire          width_adapter_007_src_endofpacket;                                                                      // width_adapter_007:out_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          width_adapter_007_src_valid;                                                                            // width_adapter_007:out_valid -> cmd_xbar_mux_005:sink1_valid
	wire          width_adapter_007_src_startofpacket;                                                                    // width_adapter_007:out_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [214:0] width_adapter_007_src_data;                                                                             // width_adapter_007:out_data -> cmd_xbar_mux_005:sink1_data
	wire          width_adapter_007_src_ready;                                                                            // cmd_xbar_mux_005:sink1_ready -> width_adapter_007:out_ready
	wire    [5:0] width_adapter_007_src_channel;                                                                          // width_adapter_007:out_channel -> cmd_xbar_mux_005:sink1_channel
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                    // rsp_xbar_demux_003:src0_endofpacket -> width_adapter_008:in_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                          // rsp_xbar_demux_003:src0_valid -> width_adapter_008:in_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                                  // rsp_xbar_demux_003:src0_startofpacket -> width_adapter_008:in_startofpacket
	wire  [214:0] rsp_xbar_demux_003_src0_data;                                                                           // rsp_xbar_demux_003:src0_data -> width_adapter_008:in_data
	wire    [5:0] rsp_xbar_demux_003_src0_channel;                                                                        // rsp_xbar_demux_003:src0_channel -> width_adapter_008:in_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                          // width_adapter_008:in_ready -> rsp_xbar_demux_003:src0_ready
	wire          width_adapter_008_src_endofpacket;                                                                      // width_adapter_008:out_endofpacket -> rsp_xbar_mux_003:sink2_endofpacket
	wire          width_adapter_008_src_valid;                                                                            // width_adapter_008:out_valid -> rsp_xbar_mux_003:sink2_valid
	wire          width_adapter_008_src_startofpacket;                                                                    // width_adapter_008:out_startofpacket -> rsp_xbar_mux_003:sink2_startofpacket
	wire  [106:0] width_adapter_008_src_data;                                                                             // width_adapter_008:out_data -> rsp_xbar_mux_003:sink2_data
	wire          width_adapter_008_src_ready;                                                                            // rsp_xbar_mux_003:sink2_ready -> width_adapter_008:out_ready
	wire    [5:0] width_adapter_008_src_channel;                                                                          // width_adapter_008:out_channel -> rsp_xbar_mux_003:sink2_channel
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                    // rsp_xbar_demux_003:src1_endofpacket -> width_adapter_009:in_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                          // rsp_xbar_demux_003:src1_valid -> width_adapter_009:in_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                                  // rsp_xbar_demux_003:src1_startofpacket -> width_adapter_009:in_startofpacket
	wire  [214:0] rsp_xbar_demux_003_src1_data;                                                                           // rsp_xbar_demux_003:src1_data -> width_adapter_009:in_data
	wire    [5:0] rsp_xbar_demux_003_src1_channel;                                                                        // rsp_xbar_demux_003:src1_channel -> width_adapter_009:in_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                          // width_adapter_009:in_ready -> rsp_xbar_demux_003:src1_ready
	wire          width_adapter_009_src_endofpacket;                                                                      // width_adapter_009:out_endofpacket -> rsp_xbar_mux_004:sink1_endofpacket
	wire          width_adapter_009_src_valid;                                                                            // width_adapter_009:out_valid -> rsp_xbar_mux_004:sink1_valid
	wire          width_adapter_009_src_startofpacket;                                                                    // width_adapter_009:out_startofpacket -> rsp_xbar_mux_004:sink1_startofpacket
	wire  [106:0] width_adapter_009_src_data;                                                                             // width_adapter_009:out_data -> rsp_xbar_mux_004:sink1_data
	wire          width_adapter_009_src_ready;                                                                            // rsp_xbar_mux_004:sink1_ready -> width_adapter_009:out_ready
	wire    [5:0] width_adapter_009_src_channel;                                                                          // width_adapter_009:out_channel -> rsp_xbar_mux_004:sink1_channel
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                    // rsp_xbar_demux_005:src0_endofpacket -> width_adapter_010:in_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                          // rsp_xbar_demux_005:src0_valid -> width_adapter_010:in_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                                  // rsp_xbar_demux_005:src0_startofpacket -> width_adapter_010:in_startofpacket
	wire  [214:0] rsp_xbar_demux_005_src0_data;                                                                           // rsp_xbar_demux_005:src0_data -> width_adapter_010:in_data
	wire    [5:0] rsp_xbar_demux_005_src0_channel;                                                                        // rsp_xbar_demux_005:src0_channel -> width_adapter_010:in_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                          // width_adapter_010:in_ready -> rsp_xbar_demux_005:src0_ready
	wire          width_adapter_010_src_endofpacket;                                                                      // width_adapter_010:out_endofpacket -> rsp_xbar_mux_003:sink4_endofpacket
	wire          width_adapter_010_src_valid;                                                                            // width_adapter_010:out_valid -> rsp_xbar_mux_003:sink4_valid
	wire          width_adapter_010_src_startofpacket;                                                                    // width_adapter_010:out_startofpacket -> rsp_xbar_mux_003:sink4_startofpacket
	wire  [106:0] width_adapter_010_src_data;                                                                             // width_adapter_010:out_data -> rsp_xbar_mux_003:sink4_data
	wire          width_adapter_010_src_ready;                                                                            // rsp_xbar_mux_003:sink4_ready -> width_adapter_010:out_ready
	wire    [5:0] width_adapter_010_src_channel;                                                                          // width_adapter_010:out_channel -> rsp_xbar_mux_003:sink4_channel
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                    // rsp_xbar_demux_005:src1_endofpacket -> width_adapter_011:in_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                          // rsp_xbar_demux_005:src1_valid -> width_adapter_011:in_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                                  // rsp_xbar_demux_005:src1_startofpacket -> width_adapter_011:in_startofpacket
	wire  [214:0] rsp_xbar_demux_005_src1_data;                                                                           // rsp_xbar_demux_005:src1_data -> width_adapter_011:in_data
	wire    [5:0] rsp_xbar_demux_005_src1_channel;                                                                        // rsp_xbar_demux_005:src1_channel -> width_adapter_011:in_channel
	wire          rsp_xbar_demux_005_src1_ready;                                                                          // width_adapter_011:in_ready -> rsp_xbar_demux_005:src1_ready
	wire          width_adapter_011_src_endofpacket;                                                                      // width_adapter_011:out_endofpacket -> rsp_xbar_mux_004:sink3_endofpacket
	wire          width_adapter_011_src_valid;                                                                            // width_adapter_011:out_valid -> rsp_xbar_mux_004:sink3_valid
	wire          width_adapter_011_src_startofpacket;                                                                    // width_adapter_011:out_startofpacket -> rsp_xbar_mux_004:sink3_startofpacket
	wire  [106:0] width_adapter_011_src_data;                                                                             // width_adapter_011:out_data -> rsp_xbar_mux_004:sink3_data
	wire          width_adapter_011_src_ready;                                                                            // rsp_xbar_mux_004:sink3_ready -> width_adapter_011:out_ready
	wire    [5:0] width_adapter_011_src_channel;                                                                          // width_adapter_011:out_channel -> rsp_xbar_mux_004:sink3_channel
	wire          cmd_xbar_demux_008_src1_ready;                                                                          // width_adapter_012:in_ready -> cmd_xbar_demux_008:src1_ready
	wire          width_adapter_012_src_endofpacket;                                                                      // width_adapter_012:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_012_src_valid;                                                                            // width_adapter_012:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_012_src_startofpacket;                                                                    // width_adapter_012:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire   [75:0] width_adapter_012_src_data;                                                                             // width_adapter_012:out_data -> burst_adapter:sink0_data
	wire          width_adapter_012_src_ready;                                                                            // burst_adapter:sink0_ready -> width_adapter_012:out_ready
	wire    [1:0] width_adapter_012_src_channel;                                                                          // width_adapter_012:out_channel -> burst_adapter:sink0_channel
	wire          id_router_019_src_endofpacket;                                                                          // id_router_019:src_endofpacket -> width_adapter_013:in_endofpacket
	wire          id_router_019_src_valid;                                                                                // id_router_019:src_valid -> width_adapter_013:in_valid
	wire          id_router_019_src_startofpacket;                                                                        // id_router_019:src_startofpacket -> width_adapter_013:in_startofpacket
	wire   [75:0] id_router_019_src_data;                                                                                 // id_router_019:src_data -> width_adapter_013:in_data
	wire    [1:0] id_router_019_src_channel;                                                                              // id_router_019:src_channel -> width_adapter_013:in_channel
	wire          id_router_019_src_ready;                                                                                // width_adapter_013:in_ready -> id_router_019:src_ready
	wire          width_adapter_013_src_endofpacket;                                                                      // width_adapter_013:out_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	wire          width_adapter_013_src_valid;                                                                            // width_adapter_013:out_valid -> rsp_xbar_demux_019:sink_valid
	wire          width_adapter_013_src_startofpacket;                                                                    // width_adapter_013:out_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	wire   [93:0] width_adapter_013_src_data;                                                                             // width_adapter_013:out_data -> rsp_xbar_demux_019:sink_data
	wire          width_adapter_013_src_ready;                                                                            // rsp_xbar_demux_019:sink_ready -> width_adapter_013:out_ready
	wire    [1:0] width_adapter_013_src_channel;                                                                          // width_adapter_013:out_channel -> rsp_xbar_demux_019:sink_channel
	wire          cmd_xbar_demux_009_src0_ready;                                                                          // width_adapter_014:in_ready -> cmd_xbar_demux_009:src0_ready
	wire          width_adapter_014_src_endofpacket;                                                                      // width_adapter_014:out_endofpacket -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          width_adapter_014_src_valid;                                                                            // width_adapter_014:out_valid -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          width_adapter_014_src_startofpacket;                                                                    // width_adapter_014:out_startofpacket -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [132:0] width_adapter_014_src_data;                                                                             // width_adapter_014:out_data -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          width_adapter_014_src_ready;                                                                            // ddr2_bot_s1_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter_014:out_ready
	wire    [0:0] width_adapter_014_src_channel;                                                                          // width_adapter_014:out_channel -> ddr2_bot_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          id_router_020_src_endofpacket;                                                                          // id_router_020:src_endofpacket -> width_adapter_015:in_endofpacket
	wire          id_router_020_src_valid;                                                                                // id_router_020:src_valid -> width_adapter_015:in_valid
	wire          id_router_020_src_startofpacket;                                                                        // id_router_020:src_startofpacket -> width_adapter_015:in_startofpacket
	wire  [132:0] id_router_020_src_data;                                                                                 // id_router_020:src_data -> width_adapter_015:in_data
	wire    [0:0] id_router_020_src_channel;                                                                              // id_router_020:src_channel -> width_adapter_015:in_channel
	wire          id_router_020_src_ready;                                                                                // width_adapter_015:in_ready -> id_router_020:src_ready
	wire          width_adapter_015_src_endofpacket;                                                                      // width_adapter_015:out_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	wire          width_adapter_015_src_valid;                                                                            // width_adapter_015:out_valid -> rsp_xbar_demux_020:sink_valid
	wire          width_adapter_015_src_startofpacket;                                                                    // width_adapter_015:out_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	wire  [204:0] width_adapter_015_src_data;                                                                             // width_adapter_015:out_data -> rsp_xbar_demux_020:sink_data
	wire          width_adapter_015_src_ready;                                                                            // rsp_xbar_demux_020:sink_ready -> width_adapter_015:out_ready
	wire    [0:0] width_adapter_015_src_channel;                                                                          // width_adapter_015:out_channel -> rsp_xbar_demux_020:sink_channel
	wire          crosser_out_endofpacket;                                                                                // crosser:out_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire          crosser_out_valid;                                                                                      // crosser:out_valid -> cmd_xbar_mux:sink0_valid
	wire          crosser_out_startofpacket;                                                                              // crosser:out_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [137:0] crosser_out_data;                                                                                       // crosser:out_data -> cmd_xbar_mux:sink0_data
	wire    [1:0] crosser_out_channel;                                                                                    // crosser:out_channel -> cmd_xbar_mux:sink0_channel
	wire          crosser_out_ready;                                                                                      // cmd_xbar_mux:sink0_ready -> crosser:out_ready
	wire          cmd_xbar_demux_src0_endofpacket;                                                                        // cmd_xbar_demux:src0_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                              // cmd_xbar_demux:src0_valid -> crosser:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                      // cmd_xbar_demux:src0_startofpacket -> crosser:in_startofpacket
	wire  [137:0] cmd_xbar_demux_src0_data;                                                                               // cmd_xbar_demux:src0_data -> crosser:in_data
	wire    [1:0] cmd_xbar_demux_src0_channel;                                                                            // cmd_xbar_demux:src0_channel -> crosser:in_channel
	wire          cmd_xbar_demux_src0_ready;                                                                              // crosser:in_ready -> cmd_xbar_demux:src0_ready
	wire          crosser_001_out_endofpacket;                                                                            // crosser_001:out_endofpacket -> width_adapter_001:in_endofpacket
	wire          crosser_001_out_valid;                                                                                  // crosser_001:out_valid -> width_adapter_001:in_valid
	wire          crosser_001_out_startofpacket;                                                                          // crosser_001:out_startofpacket -> width_adapter_001:in_startofpacket
	wire  [137:0] crosser_001_out_data;                                                                                   // crosser_001:out_data -> width_adapter_001:in_data
	wire    [1:0] crosser_001_out_channel;                                                                                // crosser_001:out_channel -> width_adapter_001:in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                        // rsp_xbar_demux:src0_endofpacket -> crosser_001:in_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                              // rsp_xbar_demux:src0_valid -> crosser_001:in_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                      // rsp_xbar_demux:src0_startofpacket -> crosser_001:in_startofpacket
	wire  [137:0] rsp_xbar_demux_src0_data;                                                                               // rsp_xbar_demux:src0_data -> crosser_001:in_data
	wire    [1:0] rsp_xbar_demux_src0_channel;                                                                            // rsp_xbar_demux:src0_channel -> crosser_001:in_channel
	wire          rsp_xbar_demux_src0_ready;                                                                              // crosser_001:in_ready -> rsp_xbar_demux:src0_ready
	wire          crosser_002_out_endofpacket;                                                                            // crosser_002:out_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire          crosser_002_out_valid;                                                                                  // crosser_002:out_valid -> cmd_xbar_mux_001:sink0_valid
	wire          crosser_002_out_startofpacket;                                                                          // crosser_002:out_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [106:0] crosser_002_out_data;                                                                                   // crosser_002:out_data -> cmd_xbar_mux_001:sink0_data
	wire    [5:0] crosser_002_out_channel;                                                                                // crosser_002:out_channel -> cmd_xbar_mux_001:sink0_channel
	wire          crosser_002_out_ready;                                                                                  // cmd_xbar_mux_001:sink0_ready -> crosser_002:out_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                    // cmd_xbar_demux_002:src0_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                          // cmd_xbar_demux_002:src0_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                                  // cmd_xbar_demux_002:src0_startofpacket -> crosser_002:in_startofpacket
	wire  [106:0] cmd_xbar_demux_002_src0_data;                                                                           // cmd_xbar_demux_002:src0_data -> crosser_002:in_data
	wire    [5:0] cmd_xbar_demux_002_src0_channel;                                                                        // cmd_xbar_demux_002:src0_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                          // crosser_002:in_ready -> cmd_xbar_demux_002:src0_ready
	wire          crosser_003_out_endofpacket;                                                                            // crosser_003:out_endofpacket -> fir_dma_read_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          crosser_003_out_valid;                                                                                  // crosser_003:out_valid -> fir_dma_read_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          crosser_003_out_startofpacket;                                                                          // crosser_003:out_startofpacket -> fir_dma_read_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [106:0] crosser_003_out_data;                                                                                   // crosser_003:out_data -> fir_dma_read_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [5:0] crosser_003_out_channel;                                                                                // crosser_003:out_channel -> fir_dma_read_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                    // rsp_xbar_demux_001:src0_endofpacket -> crosser_003:in_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                          // rsp_xbar_demux_001:src0_valid -> crosser_003:in_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                                  // rsp_xbar_demux_001:src0_startofpacket -> crosser_003:in_startofpacket
	wire  [106:0] rsp_xbar_demux_001_src0_data;                                                                           // rsp_xbar_demux_001:src0_data -> crosser_003:in_data
	wire    [5:0] rsp_xbar_demux_001_src0_channel;                                                                        // rsp_xbar_demux_001:src0_channel -> crosser_003:in_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                          // crosser_003:in_ready -> rsp_xbar_demux_001:src0_ready
	wire          crosser_004_out_endofpacket;                                                                            // crosser_004:out_endofpacket -> fir_dma_control_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_004_out_valid;                                                                                  // crosser_004:out_valid -> fir_dma_control_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_004_out_startofpacket;                                                                          // crosser_004:out_startofpacket -> fir_dma_control_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_004_out_data;                                                                                   // crosser_004:out_data -> fir_dma_control_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] crosser_004_out_channel;                                                                                // crosser_004:out_channel -> fir_dma_control_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src5_endofpacket;                                                                    // cmd_xbar_demux_007:src5_endofpacket -> crosser_004:in_endofpacket
	wire          cmd_xbar_demux_007_src5_valid;                                                                          // cmd_xbar_demux_007:src5_valid -> crosser_004:in_valid
	wire          cmd_xbar_demux_007_src5_startofpacket;                                                                  // cmd_xbar_demux_007:src5_startofpacket -> crosser_004:in_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src5_data;                                                                           // cmd_xbar_demux_007:src5_data -> crosser_004:in_data
	wire   [10:0] cmd_xbar_demux_007_src5_channel;                                                                        // cmd_xbar_demux_007:src5_channel -> crosser_004:in_channel
	wire          cmd_xbar_demux_007_src5_ready;                                                                          // crosser_004:in_ready -> cmd_xbar_demux_007:src5_ready
	wire          crosser_005_out_endofpacket;                                                                            // crosser_005:out_endofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          crosser_005_out_valid;                                                                                  // crosser_005:out_valid -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          crosser_005_out_startofpacket;                                                                          // crosser_005:out_startofpacket -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire   [82:0] crosser_005_out_data;                                                                                   // crosser_005:out_data -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire   [10:0] crosser_005_out_channel;                                                                                // crosser_005:out_channel -> pll_pll_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          cmd_xbar_demux_007_src6_endofpacket;                                                                    // cmd_xbar_demux_007:src6_endofpacket -> crosser_005:in_endofpacket
	wire          cmd_xbar_demux_007_src6_valid;                                                                          // cmd_xbar_demux_007:src6_valid -> crosser_005:in_valid
	wire          cmd_xbar_demux_007_src6_startofpacket;                                                                  // cmd_xbar_demux_007:src6_startofpacket -> crosser_005:in_startofpacket
	wire   [82:0] cmd_xbar_demux_007_src6_data;                                                                           // cmd_xbar_demux_007:src6_data -> crosser_005:in_data
	wire   [10:0] cmd_xbar_demux_007_src6_channel;                                                                        // cmd_xbar_demux_007:src6_channel -> crosser_005:in_channel
	wire          cmd_xbar_demux_007_src6_ready;                                                                          // crosser_005:in_ready -> cmd_xbar_demux_007:src6_ready
	wire          crosser_006_out_endofpacket;                                                                            // crosser_006:out_endofpacket -> rsp_xbar_mux_007:sink5_endofpacket
	wire          crosser_006_out_valid;                                                                                  // crosser_006:out_valid -> rsp_xbar_mux_007:sink5_valid
	wire          crosser_006_out_startofpacket;                                                                          // crosser_006:out_startofpacket -> rsp_xbar_mux_007:sink5_startofpacket
	wire   [82:0] crosser_006_out_data;                                                                                   // crosser_006:out_data -> rsp_xbar_mux_007:sink5_data
	wire   [10:0] crosser_006_out_channel;                                                                                // crosser_006:out_channel -> rsp_xbar_mux_007:sink5_channel
	wire          crosser_006_out_ready;                                                                                  // rsp_xbar_mux_007:sink5_ready -> crosser_006:out_ready
	wire          rsp_xbar_demux_012_src0_endofpacket;                                                                    // rsp_xbar_demux_012:src0_endofpacket -> crosser_006:in_endofpacket
	wire          rsp_xbar_demux_012_src0_valid;                                                                          // rsp_xbar_demux_012:src0_valid -> crosser_006:in_valid
	wire          rsp_xbar_demux_012_src0_startofpacket;                                                                  // rsp_xbar_demux_012:src0_startofpacket -> crosser_006:in_startofpacket
	wire   [82:0] rsp_xbar_demux_012_src0_data;                                                                           // rsp_xbar_demux_012:src0_data -> crosser_006:in_data
	wire   [10:0] rsp_xbar_demux_012_src0_channel;                                                                        // rsp_xbar_demux_012:src0_channel -> crosser_006:in_channel
	wire          rsp_xbar_demux_012_src0_ready;                                                                          // crosser_006:in_ready -> rsp_xbar_demux_012:src0_ready
	wire          crosser_007_out_endofpacket;                                                                            // crosser_007:out_endofpacket -> rsp_xbar_mux_007:sink6_endofpacket
	wire          crosser_007_out_valid;                                                                                  // crosser_007:out_valid -> rsp_xbar_mux_007:sink6_valid
	wire          crosser_007_out_startofpacket;                                                                          // crosser_007:out_startofpacket -> rsp_xbar_mux_007:sink6_startofpacket
	wire   [82:0] crosser_007_out_data;                                                                                   // crosser_007:out_data -> rsp_xbar_mux_007:sink6_data
	wire   [10:0] crosser_007_out_channel;                                                                                // crosser_007:out_channel -> rsp_xbar_mux_007:sink6_channel
	wire          crosser_007_out_ready;                                                                                  // rsp_xbar_mux_007:sink6_ready -> crosser_007:out_ready
	wire          rsp_xbar_demux_013_src0_endofpacket;                                                                    // rsp_xbar_demux_013:src0_endofpacket -> crosser_007:in_endofpacket
	wire          rsp_xbar_demux_013_src0_valid;                                                                          // rsp_xbar_demux_013:src0_valid -> crosser_007:in_valid
	wire          rsp_xbar_demux_013_src0_startofpacket;                                                                  // rsp_xbar_demux_013:src0_startofpacket -> crosser_007:in_startofpacket
	wire   [82:0] rsp_xbar_demux_013_src0_data;                                                                           // rsp_xbar_demux_013:src0_data -> crosser_007:in_data
	wire   [10:0] rsp_xbar_demux_013_src0_channel;                                                                        // rsp_xbar_demux_013:src0_channel -> crosser_007:in_channel
	wire          rsp_xbar_demux_013_src0_ready;                                                                          // crosser_007:in_ready -> rsp_xbar_demux_013:src0_ready
	wire    [5:0] limiter_cmd_valid_data;                                                                                 // limiter:cmd_src_valid -> cmd_xbar_demux_003:sink_valid
	wire    [5:0] limiter_001_cmd_valid_data;                                                                             // limiter_001:cmd_src_valid -> cmd_xbar_demux_004:sink_valid
	wire   [10:0] limiter_002_cmd_valid_data;                                                                             // limiter_002:cmd_src_valid -> cmd_xbar_demux_007:sink_valid
	wire    [1:0] limiter_003_cmd_valid_data;                                                                             // limiter_003:cmd_src_valid -> cmd_xbar_demux_008:sink_valid
	wire          irq_mapper_receiver5_irq;                                                                               // dma_0:dma_ctl_irq -> irq_mapper:receiver5_irq
	wire   [31:0] cpu_d_irq_irq;                                                                                          // irq_mapper:sender_irq -> cpu:d_irq
	wire          irq_mapper_receiver0_irq;                                                                               // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                                                          // sys_clk_timer:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver1_irq;                                                                               // irq_synchronizer_001:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                                                                      // high_res_timer:irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver2_irq;                                                                               // irq_synchronizer_002:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                                                                      // jtag_uart:av_irq -> irq_synchronizer_002:receiver_irq
	wire          irq_mapper_receiver3_irq;                                                                               // irq_synchronizer_003:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_003_receiver_irq;                                                                      // fir_dma:slave_irq -> irq_synchronizer_003:receiver_irq
	wire          irq_mapper_receiver4_irq;                                                                               // irq_synchronizer_004:sender_irq -> irq_mapper:receiver4_irq
	wire    [0:0] irq_synchronizer_004_receiver_irq;                                                                      // button_pio:irq -> irq_synchronizer_004:receiver_irq

	nios_ddr2_top ddr2_top (
		.local_address     (ddr2_top_s1_translator_avalon_anti_slave_0_address),            //                  s1.address
		.local_write_req   (ddr2_top_s1_translator_avalon_anti_slave_0_write),              //                    .write
		.local_read_req    (ddr2_top_s1_translator_avalon_anti_slave_0_read),               //                    .read
		.local_burstbegin  (ddr2_top_s1_translator_avalon_anti_slave_0_beginbursttransfer), //                    .beginbursttransfer
		.local_ready       (ddr2_top_s1_translator_avalon_anti_slave_0_waitrequest),        //                    .waitrequest_n
		.local_rdata       (ddr2_top_s1_translator_avalon_anti_slave_0_readdata),           //                    .readdata
		.local_rdata_valid (ddr2_top_s1_translator_avalon_anti_slave_0_readdatavalid),      //                    .readdatavalid
		.local_wdata       (ddr2_top_s1_translator_avalon_anti_slave_0_writedata),          //                    .writedata
		.local_be          (ddr2_top_s1_translator_avalon_anti_slave_0_byteenable),         //                    .byteenable
		.local_size        (ddr2_top_s1_translator_avalon_anti_slave_0_burstcount),         //                    .burstcount
		.local_refresh_ack (ddr2_top_external_connection_local_refresh_ack),                // external_connection.export
		.local_init_done   (ddr2_top_external_connection_local_init_done),                  //                    .export
		.reset_phy_clk_n   (ddr2_top_external_connection_reset_phy_clk_n),                  //                    .export
		.mem_odt           (ddr2_top_memory_mem_odt),                                       //              memory.mem_odt
		.mem_clk           (ddr2_top_memory_mem_clk),                                       //                    .mem_clk
		.mem_clk_n         (ddr2_top_memory_mem_clk_n),                                     //                    .mem_clk_n
		.mem_cs_n          (ddr2_top_memory_mem_cs_n),                                      //                    .mem_cs_n
		.mem_cke           (ddr2_top_memory_mem_cke),                                       //                    .mem_cke
		.mem_addr          (ddr2_top_memory_mem_addr),                                      //                    .mem_addr
		.mem_ba            (ddr2_top_memory_mem_ba),                                        //                    .mem_ba
		.mem_ras_n         (ddr2_top_memory_mem_ras_n),                                     //                    .mem_ras_n
		.mem_cas_n         (ddr2_top_memory_mem_cas_n),                                     //                    .mem_cas_n
		.mem_we_n          (ddr2_top_memory_mem_we_n),                                      //                    .mem_we_n
		.mem_dq            (ddr2_top_memory_mem_dq),                                        //                    .mem_dq
		.mem_dqs           (ddr2_top_memory_mem_dqs),                                       //                    .mem_dqs
		.mem_dm            (ddr2_top_memory_mem_dm),                                        //                    .mem_dm
		.pll_ref_clk       (clk_125),                                                       //              refclk.clk
		.soft_reset_n      (~rst_controller_reset_out_reset),                               //        soft_reset_n.reset_n
		.global_reset_n    (~rst_controller_001_reset_out_reset),                           //      global_reset_n.reset_n
		.reset_request_n   (ddr2_top_reset_request_n_reset),                                //     reset_request_n.reset_n
		.phy_clk           (sysclk_top_out_clk_clk),                                        //              sysclk.clk
		.aux_full_rate_clk (ddr2_top_auxfull_clk),                                          //             auxfull.clk
		.aux_half_rate_clk (ddr2_top_auxhalf_clk)                                           //             auxhalf.clk
	);

	nios_sys_clk_timer sys_clk_timer (
		.clk        (pll_c2_out),                                                 //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                        // reset.reset_n
		.address    (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~sys_clk_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)                               //   irq.irq
	);

	nios_high_res_timer high_res_timer (
		.clk        (pll_c2_out),                                                  //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                         // reset.reset_n
		.address    (high_res_timer_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (high_res_timer_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (high_res_timer_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (high_res_timer_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~high_res_timer_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_synchronizer_001_receiver_irq)                            //   irq.irq
	);

	nios_performance_counter performance_counter (
		.clk           (pll_c2_out),                                                                     //           clk.clk
		.reset_n       (~rst_controller_002_reset_out_reset),                                            //         reset.reset_n
		.address       (performance_counter_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.readdata      (performance_counter_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (performance_counter_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (performance_counter_control_slave_translator_avalon_anti_slave_0_writedata)      //              .writedata
	);

	nios_jtag_uart jtag_uart (
		.clk            (pll_c2_out),                                                             //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                                    //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_synchronizer_002_receiver_irq)                                       //               irq.irq
	);

	pipelined_read_burst_write_dma #(
		.DATAWIDTH                 (32),
		.BYTEENABLEWIDTH           (4),
		.ADDRESSWIDTH              (32),
		.FIFOUSEMEMORY             (1),
		.READ_FIFODEPTH            (32),
		.READ_FIFODEPTH_LOG2       (5),
		.WRITE_FIFODEPTH           (32),
		.WRITE_FIFODEPTH_LOG2      (5),
		.WRITE_MAXBURSTCOUNT       (4),
		.WRITE_MAXBURSTCOUNT_WIDTH (3)
	) fir_dma (
		.clk                       (clk),                                                       //        clock.clk
		.reset                     (rst_controller_003_reset_out_reset),                        //  clock_reset.reset
		.slave_address             (fir_dma_control_translator_avalon_anti_slave_0_address),    //      control.address
		.slave_writedata           (fir_dma_control_translator_avalon_anti_slave_0_writedata),  //             .writedata
		.slave_write               (fir_dma_control_translator_avalon_anti_slave_0_write),      //             .write
		.slave_read                (fir_dma_control_translator_avalon_anti_slave_0_read),       //             .read
		.slave_byteenable          (fir_dma_control_translator_avalon_anti_slave_0_byteenable), //             .byteenable
		.slave_readdata            (fir_dma_control_translator_avalon_anti_slave_0_readdata),   //             .readdata
		.read_master_address       (fir_dma_read_master_address),                               //  read_master.address
		.read_master_read          (fir_dma_read_master_read),                                  //             .read
		.read_master_byteenable    (fir_dma_read_master_byteenable),                            //             .byteenable
		.read_master_readdata      (fir_dma_read_master_readdata),                              //             .readdata
		.read_master_readdatavalid (fir_dma_read_master_readdatavalid),                         //             .readdatavalid
		.read_master_waitrequest   (fir_dma_read_master_waitrequest),                           //             .waitrequest
		.write_master_address      (fir_dma_write_master_address),                              // write_master.address
		.write_master_write        (fir_dma_write_master_write),                                //             .write
		.write_master_byteenable   (fir_dma_write_master_byteenable),                           //             .byteenable
		.write_master_writedata    (fir_dma_write_master_writedata),                            //             .writedata
		.write_master_waitrequest  (fir_dma_write_master_waitrequest),                          //             .waitrequest
		.write_master_burstcount   (fir_dma_write_master_burstcount),                           //             .burstcount
		.slave_irq                 (irq_synchronizer_003_receiver_irq)                          //          irq.irq
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.ADDRESS_WIDTH     (27),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) flash_ssram_pipeline_bridge (
		.clk              (pll_c0_out),                                                                  //   clk.clk
		.reset            (rst_controller_004_reset_out_reset),                                          // reset.reset
		.s0_waitrequest   (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.s0_readdatavalid (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.s0_writedata     (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.s0_address       (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_address),       //      .address
		.s0_write         (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_write),         //      .write
		.s0_read          (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_read),          //      .read
		.s0_byteenable    (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.s0_debugaccess   (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (flash_ssram_pipeline_bridge_m0_waitrequest),                                  //    m0.waitrequest
		.m0_readdata      (flash_ssram_pipeline_bridge_m0_readdata),                                     //      .readdata
		.m0_readdatavalid (flash_ssram_pipeline_bridge_m0_readdatavalid),                                //      .readdatavalid
		.m0_burstcount    (flash_ssram_pipeline_bridge_m0_burstcount),                                   //      .burstcount
		.m0_writedata     (flash_ssram_pipeline_bridge_m0_writedata),                                    //      .writedata
		.m0_address       (flash_ssram_pipeline_bridge_m0_address),                                      //      .address
		.m0_write         (flash_ssram_pipeline_bridge_m0_write),                                        //      .write
		.m0_read          (flash_ssram_pipeline_bridge_m0_read),                                         //      .read
		.m0_byteenable    (flash_ssram_pipeline_bridge_m0_byteenable),                                   //      .byteenable
		.m0_debugaccess   (flash_ssram_pipeline_bridge_m0_debugaccess)                                   //      .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (128),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (27),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) ddr2_top_clock_bridge (
		.m0_clk           (sysclk_top_out_clk_clk),                                                //   m0_clk.clk
		.m0_reset         (rst_controller_005_reset_out_reset),                                    // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                            //   s0_clk.clk
		.s0_reset         (rst_controller_004_reset_out_reset),                                    // s0_reset.reset
		.s0_waitrequest   (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (ddr2_top_clock_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (ddr2_top_clock_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (ddr2_top_clock_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (ddr2_top_clock_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (ddr2_top_clock_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (ddr2_top_clock_bridge_m0_address),                                      //         .address
		.m0_write         (ddr2_top_clock_bridge_m0_write),                                        //         .write
		.m0_read          (ddr2_top_clock_bridge_m0_read),                                         //         .read
		.m0_byteenable    (ddr2_top_clock_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (ddr2_top_clock_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (16),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) slow_peripheral_bridge (
		.m0_clk           (pll_c2_out),                                                             //   m0_clk.clk
		.m0_reset         (rst_controller_002_reset_out_reset),                                     // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                             //   s0_clk.clk
		.s0_reset         (rst_controller_004_reset_out_reset),                                     // s0_reset.reset
		.s0_waitrequest   (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (slow_peripheral_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (slow_peripheral_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (slow_peripheral_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (slow_peripheral_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (slow_peripheral_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (slow_peripheral_bridge_m0_address),                                      //         .address
		.m0_write         (slow_peripheral_bridge_m0_write),                                        //         .write
		.m0_read          (slow_peripheral_bridge_m0_read),                                         //         .read
		.m0_byteenable    (slow_peripheral_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (slow_peripheral_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	nios_sysid sysid (
		.clock    (pll_c2_out),                                                  //           clk.clk
		.reset_n  (~rst_controller_002_reset_out_reset),                         //         reset.reset_n
		.readdata (sysid_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	nios_flash_ssram_tristate_bridge_bridge_0 flash_ssram_tristate_bridge_bridge_0 (
		.clk                                        (pll_c0_out),                                                                          //   clk.clk
		.reset                                      (rst_controller_004_reset_out_reset),                                                  // reset.reset
		.request                                    (flash_ssram_tristate_bridge_pinsharer_0_tcm_request),                                 //   tcs.request
		.grant                                      (flash_ssram_tristate_bridge_pinsharer_0_tcm_grant),                                   //      .grant
		.tcs_read_n_to_the_ext_flash                (flash_ssram_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out),             //      .read_n_to_the_ext_flash_out
		.tcs_select_n_to_the_ext_flash              (flash_ssram_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out),           //      .select_n_to_the_ext_flash_out
		.tcs_flash_ssram_tristate_bridge_address    (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_address_out), //      .flash_ssram_tristate_bridge_address_out
		.tcs_bwe_n_to_the_ssram                     (flash_ssram_tristate_bridge_pinsharer_0_tcm_bwe_n_to_the_ssram_out),                  //      .bwe_n_to_the_ssram_out
		.tcs_reset_n_to_the_ssram                   (flash_ssram_tristate_bridge_pinsharer_0_tcm_reset_n_to_the_ssram_out),                //      .reset_n_to_the_ssram_out
		.tcs_chipenable1_n_to_the_ssram             (flash_ssram_tristate_bridge_pinsharer_0_tcm_chipenable1_n_to_the_ssram_out),          //      .chipenable1_n_to_the_ssram_out
		.tcs_bw_n_to_the_ssram                      (flash_ssram_tristate_bridge_pinsharer_0_tcm_bw_n_to_the_ssram_out),                   //      .bw_n_to_the_ssram_out
		.tcs_outputenable_n_to_the_ssram            (flash_ssram_tristate_bridge_pinsharer_0_tcm_outputenable_n_to_the_ssram_out),         //      .outputenable_n_to_the_ssram_out
		.tcs_flash_ssram_tristate_bridge_data       (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_out),    //      .flash_ssram_tristate_bridge_data_out
		.tcs_flash_ssram_tristate_bridge_data_outen (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_outen),  //      .flash_ssram_tristate_bridge_data_outen
		.tcs_flash_ssram_tristate_bridge_data_in    (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_in),     //      .flash_ssram_tristate_bridge_data_in
		.tcs_adsc_n_to_the_ssram                    (flash_ssram_tristate_bridge_pinsharer_0_tcm_adsc_n_to_the_ssram_out),                 //      .adsc_n_to_the_ssram_out
		.tcs_address_to_the_ssram                   (flash_ssram_tristate_bridge_pinsharer_0_tcm_address_to_the_ssram_out),                //      .address_to_the_ssram_out
		.tcs_write_n_to_the_ext_flash               (flash_ssram_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out),            //      .write_n_to_the_ext_flash_out
		.read_n_to_the_ext_flash                    (read_n_to_the_ext_flash),                                                             //   out.read_n_to_the_ext_flash
		.select_n_to_the_ext_flash                  (select_n_to_the_ext_flash),                                                           //      .select_n_to_the_ext_flash
		.flash_ssram_tristate_bridge_address        (flash_ssram_tristate_bridge_address),                                                 //      .flash_ssram_tristate_bridge_address
		.bwe_n_to_the_ssram                         (bwe_n_to_the_ssram),                                                                  //      .bwe_n_to_the_ssram
		.reset_n_to_the_ssram                       (reset_n_to_the_ssram),                                                                //      .reset_n_to_the_ssram
		.chipenable1_n_to_the_ssram                 (chipenable1_n_to_the_ssram),                                                          //      .chipenable1_n_to_the_ssram
		.bw_n_to_the_ssram                          (bw_n_to_the_ssram),                                                                   //      .bw_n_to_the_ssram
		.outputenable_n_to_the_ssram                (outputenable_n_to_the_ssram),                                                         //      .outputenable_n_to_the_ssram
		.flash_ssram_tristate_bridge_data           (flash_ssram_tristate_bridge_data),                                                    //      .flash_ssram_tristate_bridge_data
		.adsc_n_to_the_ssram                        (adsc_n_to_the_ssram),                                                                 //      .adsc_n_to_the_ssram
		.address_to_the_ssram                       (address_to_the_ssram),                                                                //      .address_to_the_ssram
		.write_n_to_the_ext_flash                   (write_n_to_the_ext_flash)                                                             //      .write_n_to_the_ext_flash
	);

	nios_flash_ssram_tristate_bridge_pinSharer_0 flash_ssram_tristate_bridge_pinsharer_0 (
		.clk_clk                                (pll_c0_out),                                                                          //   clk.clk
		.reset_reset                            (rst_controller_004_reset_out_reset),                                                  // reset.reset
		.request                                (flash_ssram_tristate_bridge_pinsharer_0_tcm_request),                                 //   tcm.request
		.grant                                  (flash_ssram_tristate_bridge_pinsharer_0_tcm_grant),                                   //      .grant
		.flash_ssram_tristate_bridge_address    (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_address_out), //      .flash_ssram_tristate_bridge_address_out
		.read_n_to_the_ext_flash                (flash_ssram_tristate_bridge_pinsharer_0_tcm_read_n_to_the_ext_flash_out),             //      .read_n_to_the_ext_flash_out
		.write_n_to_the_ext_flash               (flash_ssram_tristate_bridge_pinsharer_0_tcm_write_n_to_the_ext_flash_out),            //      .write_n_to_the_ext_flash_out
		.select_n_to_the_ext_flash              (flash_ssram_tristate_bridge_pinsharer_0_tcm_select_n_to_the_ext_flash_out),           //      .select_n_to_the_ext_flash_out
		.chipenable1_n_to_the_ssram             (flash_ssram_tristate_bridge_pinsharer_0_tcm_chipenable1_n_to_the_ssram_out),          //      .chipenable1_n_to_the_ssram_out
		.bw_n_to_the_ssram                      (flash_ssram_tristate_bridge_pinsharer_0_tcm_bw_n_to_the_ssram_out),                   //      .bw_n_to_the_ssram_out
		.outputenable_n_to_the_ssram            (flash_ssram_tristate_bridge_pinsharer_0_tcm_outputenable_n_to_the_ssram_out),         //      .outputenable_n_to_the_ssram_out
		.bwe_n_to_the_ssram                     (flash_ssram_tristate_bridge_pinsharer_0_tcm_bwe_n_to_the_ssram_out),                  //      .bwe_n_to_the_ssram_out
		.flash_ssram_tristate_bridge_data       (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_out),    //      .flash_ssram_tristate_bridge_data_out
		.flash_ssram_tristate_bridge_data_in    (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_in),     //      .flash_ssram_tristate_bridge_data_in
		.flash_ssram_tristate_bridge_data_outen (flash_ssram_tristate_bridge_pinsharer_0_tcm_flash_ssram_tristate_bridge_data_outen),  //      .flash_ssram_tristate_bridge_data_outen
		.address_to_the_ssram                   (flash_ssram_tristate_bridge_pinsharer_0_tcm_address_to_the_ssram_out),                //      .address_to_the_ssram_out
		.reset_n_to_the_ssram                   (flash_ssram_tristate_bridge_pinsharer_0_tcm_reset_n_to_the_ssram_out),                //      .reset_n_to_the_ssram_out
		.adsc_n_to_the_ssram                    (flash_ssram_tristate_bridge_pinsharer_0_tcm_adsc_n_to_the_ssram_out),                 //      .adsc_n_to_the_ssram_out
		.tcs0_request                           (ssram_tcm_request),                                                                   //  tcs0.request
		.tcs0_grant                             (ssram_tcm_grant),                                                                     //      .grant
		.tcs0_chipselect_n_out                  (ssram_tcm_chipselect_n_out),                                                          //      .chipselect_n_out
		.tcs0_byteenable_n_out                  (ssram_tcm_byteenable_n_out),                                                          //      .byteenable_n_out
		.tcs0_outputenable_n_out                (ssram_tcm_outputenable_n_out),                                                        //      .outputenable_n_out
		.tcs0_write_n_out                       (ssram_tcm_write_n_out),                                                               //      .write_n_out
		.tcs0_data_out                          (ssram_tcm_data_out),                                                                  //      .data_out
		.tcs0_data_in                           (ssram_tcm_data_in),                                                                   //      .data_in
		.tcs0_data_outen                        (ssram_tcm_data_outen),                                                                //      .data_outen
		.tcs0_address_out                       (ssram_tcm_address_out),                                                               //      .address_out
		.tcs0_reset_n_out                       (ssram_tcm_reset_n_out),                                                               //      .reset_n_out
		.tcs0_begintransfer_n_out               (ssram_tcm_begintransfer_n_out),                                                       //      .begintransfer_n_out
		.tcs1_request                           (ext_flash_tcm_request),                                                               //  tcs1.request
		.tcs1_grant                             (ext_flash_tcm_grant),                                                                 //      .grant
		.tcs1_address_out                       (ext_flash_tcm_address_out),                                                           //      .address_out
		.tcs1_read_n_out                        (ext_flash_tcm_read_n_out),                                                            //      .read_n_out
		.tcs1_write_n_out                       (ext_flash_tcm_write_n_out),                                                           //      .write_n_out
		.tcs1_data_out                          (ext_flash_tcm_data_out),                                                              //      .data_out
		.tcs1_data_in                           (ext_flash_tcm_data_in),                                                               //      .data_in
		.tcs1_data_outen                        (ext_flash_tcm_data_outen),                                                            //      .data_outen
		.tcs1_chipselect_n_out                  (ext_flash_tcm_chipselect_n_out)                                                       //      .chipselect_n_out
	);

	nios_ssram #(
		.TCM_ADDRESS_W                  (20),
		.TCM_DATA_W                     (32),
		.TCM_BYTEENABLE_W               (4),
		.TCM_READ_WAIT                  (0),
		.TCM_WRITE_WAIT                 (0),
		.TCM_SETUP_WAIT                 (0),
		.TCM_DATA_HOLD                  (0),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (1),
		.TCM_READLATENCY                (4),
		.TCM_SYMBOLS_PER_WORD           (4),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (1),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (1),
		.CHIPSELECT_THROUGH_READLATENCY (1)
	) ssram (
		.clk_clk                 (pll_c0_out),                                             //   clk.clk
		.reset_reset             (rst_controller_004_reset_out_reset),                     // reset.reset
		.uas_address             (ssram_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount          (ssram_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read                (ssram_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write               (ssram_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest         (ssram_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid       (ssram_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable          (ssram_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata            (ssram_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata           (ssram_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock                (ssram_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess         (ssram_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out         (ssram_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_begintransfer_n_out (ssram_tcm_begintransfer_n_out),                          //      .begintransfer_n_out
		.tcm_chipselect_n_out    (ssram_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_outputenable_n_out  (ssram_tcm_outputenable_n_out),                           //      .outputenable_n_out
		.tcm_reset_n_out         (ssram_tcm_reset_n_out),                                  //      .reset_n_out
		.tcm_request             (ssram_tcm_request),                                      //      .request
		.tcm_grant               (ssram_tcm_grant),                                        //      .grant
		.tcm_address_out         (ssram_tcm_address_out),                                  //      .address_out
		.tcm_byteenable_n_out    (ssram_tcm_byteenable_n_out),                             //      .byteenable_n_out
		.tcm_data_out            (ssram_tcm_data_out),                                     //      .data_out
		.tcm_data_outen          (ssram_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in             (ssram_tcm_data_in)                                       //      .data_in
	);

	nios_ext_flash #(
		.TCM_ADDRESS_W                  (26),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (40),
		.TCM_WRITE_WAIT                 (40),
		.TCM_SETUP_WAIT                 (80),
		.TCM_DATA_HOLD                  (20),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) ext_flash (
		.clk_clk              (pll_c0_out),                                                 //   clk.clk
		.reset_reset          (rst_controller_004_reset_out_reset),                         // reset.reset
		.uas_address          (ext_flash_uas_translator_avalon_anti_slave_0_address),       //   uas.address
		.uas_burstcount       (ext_flash_uas_translator_avalon_anti_slave_0_burstcount),    //      .burstcount
		.uas_read             (ext_flash_uas_translator_avalon_anti_slave_0_read),          //      .read
		.uas_write            (ext_flash_uas_translator_avalon_anti_slave_0_write),         //      .write
		.uas_waitrequest      (ext_flash_uas_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.uas_byteenable       (ext_flash_uas_translator_avalon_anti_slave_0_byteenable),    //      .byteenable
		.uas_readdata         (ext_flash_uas_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.uas_writedata        (ext_flash_uas_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.uas_lock             (ext_flash_uas_translator_avalon_anti_slave_0_lock),          //      .lock
		.uas_debugaccess      (ext_flash_uas_translator_avalon_anti_slave_0_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (ext_flash_tcm_write_n_out),                                  //   tcm.write_n_out
		.tcm_read_n_out       (ext_flash_tcm_read_n_out),                                   //      .read_n_out
		.tcm_chipselect_n_out (ext_flash_tcm_chipselect_n_out),                             //      .chipselect_n_out
		.tcm_request          (ext_flash_tcm_request),                                      //      .request
		.tcm_grant            (ext_flash_tcm_grant),                                        //      .grant
		.tcm_address_out      (ext_flash_tcm_address_out),                                  //      .address_out
		.tcm_data_out         (ext_flash_tcm_data_out),                                     //      .data_out
		.tcm_data_outen       (ext_flash_tcm_data_outen),                                   //      .data_outen
		.tcm_data_in          (ext_flash_tcm_data_in)                                       //      .data_in
	);

	nios_cpu cpu (
		.clk                                   (pll_c0_out),                                                       //                       clk.clk
		.reset_n                               (~rst_controller_004_reset_out_reset),                              //                   reset_n.reset_n
		.d_address                             (cpu_data_master_address),                                          //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                                       //                          .byteenable
		.d_read                                (cpu_data_master_read),                                             //                          .read
		.d_readdata                            (cpu_data_master_readdata),                                         //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                                      //                          .waitrequest
		.d_write                               (cpu_data_master_write),                                            //                          .write
		.d_writedata                           (cpu_data_master_writedata),                                        //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                                    //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                                      //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                                   //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                                      //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                                  //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                               //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                             //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                                    //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                                //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),        //                          .read
		.jtag_debug_module_readdata            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),       //                          .write
		.jtag_debug_module_writedata           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                                  // custom_instruction_master.readra
	);

	nios_pll pll (
		.clk       (clk),                                                    //       inclk_interface.clk
		.reset     (rst_controller_003_reset_out_reset),                     // inclk_interface_reset.reset
		.read      (pll_pll_slave_translator_avalon_anti_slave_0_read),      //             pll_slave.read
		.write     (pll_pll_slave_translator_avalon_anti_slave_0_write),     //                      .write
		.address   (pll_pll_slave_translator_avalon_anti_slave_0_address),   //                      .address
		.readdata  (pll_pll_slave_translator_avalon_anti_slave_0_readdata),  //                      .readdata
		.writedata (pll_pll_slave_translator_avalon_anti_slave_0_writedata), //                      .writedata
		.c0        (pll_c0_out),                                             //                    c0.clk
		.c2        (pll_c2_out),                                             //                    c2.clk
		.areset    (),                                                       //        areset_conduit.export
		.locked    (),                                                       //        locked_conduit.export
		.phasedone ()                                                        //     phasedone_conduit.export
	);

	nios_button_pio button_pio (
		.clk        (pll_c2_out),                                              //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                     //               reset.reset_n
		.address    (button_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),                   // external_connection.export
		.irq        (irq_synchronizer_004_receiver_irq)                        //                 irq.irq
	);

	nios_led_pio led_pio (
		.clk        (pll_c2_out),                                           //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                  //               reset.reset_n
		.address    (led_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)                    // external_connection.export
	);

	nios_lcd_display lcd_display (
		.reset_n       (~rst_controller_002_reset_out_reset),                                    //         reset.reset_n
		.clk           (pll_c2_out),                                                             //           clk.clk
		.begintransfer (lcd_display_control_slave_translator_avalon_anti_slave_0_begintransfer), // control_slave.begintransfer
		.read          (lcd_display_control_slave_translator_avalon_anti_slave_0_read),          //              .read
		.write         (lcd_display_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.readdata      (lcd_display_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.writedata     (lcd_display_control_slave_translator_avalon_anti_slave_0_writedata),     //              .writedata
		.address       (lcd_display_control_slave_translator_avalon_anti_slave_0_address),       //              .address
		.LCD_RS        (lcd_display_external_RS),                                                //      external.export
		.LCD_RW        (lcd_display_external_RW),                                                //              .export
		.LCD_data      (lcd_display_external_data),                                              //              .export
		.LCD_E         (lcd_display_external_E)                                                  //              .export
	);

	nios_seven_seg_pio seven_seg_pio (
		.clk        (pll_c2_out),                                                 //                 clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),                        //               reset.reset_n
		.address    (seven_seg_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~seven_seg_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (seven_seg_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (seven_seg_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (seven_seg_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (seven_seg_pio_external_connection_export)                    // external_connection.export
	);

	nios_ddr2_top ddr2_bot (
		.local_address     (ddr2_bot_s1_translator_avalon_anti_slave_0_address),            //                  s1.address
		.local_write_req   (ddr2_bot_s1_translator_avalon_anti_slave_0_write),              //                    .write
		.local_read_req    (ddr2_bot_s1_translator_avalon_anti_slave_0_read),               //                    .read
		.local_burstbegin  (ddr2_bot_s1_translator_avalon_anti_slave_0_beginbursttransfer), //                    .beginbursttransfer
		.local_ready       (ddr2_bot_s1_translator_avalon_anti_slave_0_waitrequest),        //                    .waitrequest_n
		.local_rdata       (ddr2_bot_s1_translator_avalon_anti_slave_0_readdata),           //                    .readdata
		.local_rdata_valid (ddr2_bot_s1_translator_avalon_anti_slave_0_readdatavalid),      //                    .readdatavalid
		.local_wdata       (ddr2_bot_s1_translator_avalon_anti_slave_0_writedata),          //                    .writedata
		.local_be          (ddr2_bot_s1_translator_avalon_anti_slave_0_byteenable),         //                    .byteenable
		.local_size        (ddr2_bot_s1_translator_avalon_anti_slave_0_burstcount),         //                    .burstcount
		.local_refresh_ack (ddr2_bot_external_connection_local_refresh_ack),                // external_connection.export
		.local_init_done   (ddr2_bot_external_connection_local_init_done),                  //                    .export
		.reset_phy_clk_n   (ddr2_bot_external_connection_reset_phy_clk_n),                  //                    .export
		.mem_odt           (ddr2_bot_memory_mem_odt),                                       //              memory.mem_odt
		.mem_clk           (ddr2_bot_memory_mem_clk),                                       //                    .mem_clk
		.mem_clk_n         (ddr2_bot_memory_mem_clk_n),                                     //                    .mem_clk_n
		.mem_cs_n          (ddr2_bot_memory_mem_cs_n),                                      //                    .mem_cs_n
		.mem_cke           (ddr2_bot_memory_mem_cke),                                       //                    .mem_cke
		.mem_addr          (ddr2_bot_memory_mem_addr),                                      //                    .mem_addr
		.mem_ba            (ddr2_bot_memory_mem_ba),                                        //                    .mem_ba
		.mem_ras_n         (ddr2_bot_memory_mem_ras_n),                                     //                    .mem_ras_n
		.mem_cas_n         (ddr2_bot_memory_mem_cas_n),                                     //                    .mem_cas_n
		.mem_we_n          (ddr2_bot_memory_mem_we_n),                                      //                    .mem_we_n
		.mem_dq            (ddr2_bot_memory_mem_dq),                                        //                    .mem_dq
		.mem_dqs           (ddr2_bot_memory_mem_dqs),                                       //                    .mem_dqs
		.mem_dm            (ddr2_bot_memory_mem_dm),                                        //                    .mem_dm
		.pll_ref_clk       (clk_125),                                                       //              refclk.clk
		.soft_reset_n      (~rst_controller_reset_out_reset),                               //        soft_reset_n.reset_n
		.global_reset_n    (~rst_controller_001_reset_out_reset),                           //      global_reset_n.reset_n
		.reset_request_n   (ddr2_bot_reset_request_n_reset),                                //     reset_request_n.reset_n
		.phy_clk           (sysclk_bot_out_clk_clk),                                        //              sysclk.clk
		.aux_full_rate_clk (),                                                              //             auxfull.clk
		.aux_half_rate_clk ()                                                               //             auxhalf.clk
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (128),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (27),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) ddr2_bot_clock_bridge (
		.m0_clk           (sysclk_bot_out_clk_clk),                                                //   m0_clk.clk
		.m0_reset         (rst_controller_006_reset_out_reset),                                    // m0_reset.reset
		.s0_clk           (pll_c0_out),                                                            //   s0_clk.clk
		.s0_reset         (rst_controller_004_reset_out_reset),                                    // s0_reset.reset
		.s0_waitrequest   (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),      //         .readdata
		.s0_readdatavalid (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),    //         .burstcount
		.s0_writedata     (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),     //         .writedata
		.s0_address       (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_address),       //         .address
		.s0_write         (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_write),         //         .write
		.s0_read          (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_read),          //         .read
		.s0_byteenable    (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),    //         .byteenable
		.s0_debugaccess   (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (ddr2_bot_clock_bridge_m0_waitrequest),                                  //       m0.waitrequest
		.m0_readdata      (ddr2_bot_clock_bridge_m0_readdata),                                     //         .readdata
		.m0_readdatavalid (ddr2_bot_clock_bridge_m0_readdatavalid),                                //         .readdatavalid
		.m0_burstcount    (ddr2_bot_clock_bridge_m0_burstcount),                                   //         .burstcount
		.m0_writedata     (ddr2_bot_clock_bridge_m0_writedata),                                    //         .writedata
		.m0_address       (ddr2_bot_clock_bridge_m0_address),                                      //         .address
		.m0_write         (ddr2_bot_clock_bridge_m0_write),                                        //         .write
		.m0_read          (ddr2_bot_clock_bridge_m0_read),                                         //         .read
		.m0_byteenable    (ddr2_bot_clock_bridge_m0_byteenable),                                   //         .byteenable
		.m0_debugaccess   (ddr2_bot_clock_bridge_m0_debugaccess)                                   //         .debugaccess
	);

	nios_dma_0 dma_0 (
		.clk                (pll_c0_out),                                                         //                clk.clk
		.system_reset_n     (~rst_controller_004_reset_out_reset),                                //              reset.reset_n
		.dma_ctl_address    (dma_0_control_port_slave_translator_avalon_anti_slave_0_address),    // control_port_slave.address
		.dma_ctl_chipselect (dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect), //                   .chipselect
		.dma_ctl_readdata   (dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata),   //                   .readdata
		.dma_ctl_write_n    (~dma_0_control_port_slave_translator_avalon_anti_slave_0_write),     //                   .write_n
		.dma_ctl_writedata  (dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata),  //                   .writedata
		.dma_ctl_irq        (irq_mapper_receiver5_irq),                                           //                irq.irq
		.read_address       (dma_0_read_master_address),                                          //        read_master.address
		.read_chipselect    (dma_0_read_master_chipselect),                                       //                   .chipselect
		.read_read_n        (dma_0_read_master_read),                                             //                   .read_n
		.read_readdata      (dma_0_read_master_readdata),                                         //                   .readdata
		.read_readdatavalid (dma_0_read_master_readdatavalid),                                    //                   .readdatavalid
		.read_waitrequest   (dma_0_read_master_waitrequest),                                      //                   .waitrequest
		.write_address      (dma_0_write_master_address),                                         //       write_master.address
		.write_chipselect   (dma_0_write_master_chipselect),                                      //                   .chipselect
		.write_waitrequest  (dma_0_write_master_waitrequest),                                     //                   .waitrequest
		.write_write_n      (dma_0_write_master_write),                                           //                   .write_n
		.write_writedata    (dma_0_write_master_writedata),                                       //                   .writedata
		.write_byteenable   (dma_0_write_master_byteenable)                                       //                   .byteenable
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (3),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (5),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) fir_dma_write_master_translator (
		.clk                      (clk),                                                                     //                       clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                      //                     reset.reset
		.uav_address              (fir_dma_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (fir_dma_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (fir_dma_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (fir_dma_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (fir_dma_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (fir_dma_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (fir_dma_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (fir_dma_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (fir_dma_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (fir_dma_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (fir_dma_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (fir_dma_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (fir_dma_write_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (fir_dma_write_master_burstcount),                                         //                          .burstcount
		.av_byteenable            (fir_dma_write_master_byteenable),                                         //                          .byteenable
		.av_write                 (fir_dma_write_master_write),                                              //                          .write
		.av_writedata             (fir_dma_write_master_writedata),                                          //                          .writedata
		.av_beginbursttransfer    (1'b0),                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                    //               (terminated)
		.av_read                  (1'b0),                                                                    //               (terminated)
		.av_readdata              (),                                                                        //               (terminated)
		.av_readdatavalid         (),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                    //               (terminated)
		.av_debugaccess           (1'b0),                                                                    //               (terminated)
		.uav_clken                (),                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                   //               (terminated)
		.av_response              (),                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                         //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (128),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (16),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (5),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (16),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) ddr2_top_clock_bridge_m0_translator (
		.clk                      (sysclk_top_out_clk_clk),                                                      //                       clk.clk
		.reset                    (rst_controller_005_reset_out_reset),                                          //                     reset.reset
		.uav_address              (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (ddr2_top_clock_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (ddr2_top_clock_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (ddr2_top_clock_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (ddr2_top_clock_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read                  (ddr2_top_clock_bridge_m0_read),                                               //                          .read
		.av_readdata              (ddr2_top_clock_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (ddr2_top_clock_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (ddr2_top_clock_bridge_m0_write),                                              //                          .write
		.av_writedata             (ddr2_top_clock_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (ddr2_top_clock_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (6),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_top_s1_translator (
		.clk                      (sysclk_top_out_clk_clk),                                                 //                      clk.clk
		.reset                    (~ddr2_top_reset_request_n_reset),                                        //                    reset.reset
		.uav_address              (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_top_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_top_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ddr2_top_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ddr2_top_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_top_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer    (ddr2_top_s1_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount            (ddr2_top_s1_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ddr2_top_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ddr2_top_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (~ddr2_top_s1_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) fir_dma_read_master_translator (
		.clk                      (clk),                                                                    //                       clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                     //                     reset.reset
		.uav_address              (fir_dma_read_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (fir_dma_read_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (fir_dma_read_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (fir_dma_read_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (fir_dma_read_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (fir_dma_read_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (fir_dma_read_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (fir_dma_read_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (fir_dma_read_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (fir_dma_read_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (fir_dma_read_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (fir_dma_read_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (fir_dma_read_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (fir_dma_read_master_byteenable),                                         //                          .byteenable
		.av_read                  (fir_dma_read_master_read),                                               //                          .read
		.av_readdata              (fir_dma_read_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (fir_dma_read_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                   //               (terminated)
		.av_begintransfer         (1'b0),                                                                   //               (terminated)
		.av_chipselect            (1'b0),                                                                   //               (terminated)
		.av_write                 (1'b0),                                                                   //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                   //               (terminated)
		.av_lock                  (1'b0),                                                                   //               (terminated)
		.av_debugaccess           (1'b0),                                                                   //               (terminated)
		.uav_clken                (),                                                                       //               (terminated)
		.av_clken                 (1'b1),                                                                   //               (terminated)
		.uav_response             (2'b00),                                                                  //               (terminated)
		.av_response              (),                                                                       //               (terminated)
		.uav_writeresponserequest (),                                                                       //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                   //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                   //               (terminated)
		.av_writeresponsevalid    ()                                                                        //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_data_master_translator (
		.clk                      (pll_c0_out),                                                         //                       clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                 //                     reset.reset
		.uav_address              (cpu_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (cpu_data_master_byteenable),                                         //                          .byteenable
		.av_read                  (cpu_data_master_read),                                               //                          .read
		.av_readdata              (cpu_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (cpu_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (cpu_data_master_write),                                              //                          .write
		.av_writedata             (cpu_data_master_writedata),                                          //                          .writedata
		.av_debugaccess           (cpu_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount            (1'b1),                                                               //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                               //               (terminated)
		.av_begintransfer         (1'b0),                                                               //               (terminated)
		.av_chipselect            (1'b0),                                                               //               (terminated)
		.av_lock                  (1'b0),                                                               //               (terminated)
		.uav_clken                (),                                                                   //               (terminated)
		.av_clken                 (1'b1),                                                               //               (terminated)
		.uav_response             (2'b00),                                                              //               (terminated)
		.av_response              (),                                                                   //               (terminated)
		.uav_writeresponserequest (),                                                                   //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                               //               (terminated)
		.av_writeresponserequest  (1'b0),                                                               //               (terminated)
		.av_writeresponsevalid    ()                                                                    //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) cpu_instruction_master_translator (
		.clk                      (pll_c0_out),                                                                //                       clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                        //                     reset.reset
		.uav_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (cpu_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (cpu_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read                  (cpu_instruction_master_read),                                               //                          .read
		.av_readdata              (cpu_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (cpu_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                      //               (terminated)
		.av_byteenable            (4'b1111),                                                                   //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                      //               (terminated)
		.av_begintransfer         (1'b0),                                                                      //               (terminated)
		.av_chipselect            (1'b0),                                                                      //               (terminated)
		.av_write                 (1'b0),                                                                      //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                      //               (terminated)
		.av_lock                  (1'b0),                                                                      //               (terminated)
		.av_debugaccess           (1'b0),                                                                      //               (terminated)
		.uav_clken                (),                                                                          //               (terminated)
		.av_clken                 (1'b1),                                                                      //               (terminated)
		.uav_response             (2'b00),                                                                     //               (terminated)
		.av_response              (),                                                                          //               (terminated)
		.uav_writeresponserequest (),                                                                          //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                      //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                      //               (terminated)
		.av_writeresponsevalid    ()                                                                           //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (30),
		.AV_DATA_W                   (128),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (16),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (5),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (16),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_0_read_master_translator (
		.clk                      (pll_c0_out),                                                                                                                            //                       clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                                                                                    //                     reset.reset
		.uav_address              (dma_0_read_master_translator_avalon_universal_master_0_address),                                                                        // avalon_universal_master_0.address
		.uav_burstcount           (dma_0_read_master_translator_avalon_universal_master_0_burstcount),                                                                     //                          .burstcount
		.uav_read                 (dma_0_read_master_translator_avalon_universal_master_0_read),                                                                           //                          .read
		.uav_write                (dma_0_read_master_translator_avalon_universal_master_0_write),                                                                          //                          .write
		.uav_waitrequest          (dma_0_read_master_translator_avalon_universal_master_0_waitrequest),                                                                    //                          .waitrequest
		.uav_readdatavalid        (dma_0_read_master_translator_avalon_universal_master_0_readdatavalid),                                                                  //                          .readdatavalid
		.uav_byteenable           (dma_0_read_master_translator_avalon_universal_master_0_byteenable),                                                                     //                          .byteenable
		.uav_readdata             (dma_0_read_master_translator_avalon_universal_master_0_readdata),                                                                       //                          .readdata
		.uav_writedata            (dma_0_read_master_translator_avalon_universal_master_0_writedata),                                                                      //                          .writedata
		.uav_lock                 (dma_0_read_master_translator_avalon_universal_master_0_lock),                                                                           //                          .lock
		.uav_debugaccess          (dma_0_read_master_translator_avalon_universal_master_0_debugaccess),                                                                    //                          .debugaccess
		.av_address               (dma_0_read_master_address),                                                                                                             //      avalon_anti_master_0.address
		.av_waitrequest           (dma_0_read_master_waitrequest),                                                                                                         //                          .waitrequest
		.av_chipselect            (dma_0_read_master_chipselect),                                                                                                          //                          .chipselect
		.av_read                  (~dma_0_read_master_read),                                                                                                               //                          .read
		.av_readdata              (dma_0_read_master_readdata),                                                                                                            //                          .readdata
		.av_readdatavalid         (dma_0_read_master_readdatavalid),                                                                                                       //                          .readdatavalid
		.av_burstcount            (1'b1),                                                                                                                                  //               (terminated)
		.av_byteenable            (16'b1111111111111111),                                                                                                                  //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                                                                                  //               (terminated)
		.av_write                 (1'b0),                                                                                                                                  //               (terminated)
		.av_writedata             (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //               (terminated)
		.av_lock                  (1'b0),                                                                                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                                                                                  //               (terminated)
		.uav_clken                (),                                                                                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                                                                                 //               (terminated)
		.av_response              (),                                                                                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                                                                                       //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (29),
		.AV_DATA_W                   (128),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (16),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (5),
		.USE_READ                    (0),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (1),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (0),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (16),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) dma_0_write_master_translator (
		.clk                      (pll_c0_out),                                                            //                       clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                    //                     reset.reset
		.uav_address              (dma_0_write_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (dma_0_write_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (dma_0_write_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (dma_0_write_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (dma_0_write_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (dma_0_write_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (dma_0_write_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (dma_0_write_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (dma_0_write_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (dma_0_write_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (dma_0_write_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (dma_0_write_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (dma_0_write_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (dma_0_write_master_byteenable),                                         //                          .byteenable
		.av_chipselect            (dma_0_write_master_chipselect),                                         //                          .chipselect
		.av_write                 (~dma_0_write_master_write),                                             //                          .write
		.av_writedata             (dma_0_write_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                  //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                  //               (terminated)
		.av_begintransfer         (1'b0),                                                                  //               (terminated)
		.av_read                  (1'b0),                                                                  //               (terminated)
		.av_readdata              (),                                                                      //               (terminated)
		.av_readdatavalid         (),                                                                      //               (terminated)
		.av_lock                  (1'b0),                                                                  //               (terminated)
		.av_debugaccess           (1'b0),                                                                  //               (terminated)
		.uav_clken                (),                                                                      //               (terminated)
		.av_clken                 (1'b1),                                                                  //               (terminated)
		.uav_response             (2'b00),                                                                 //               (terminated)
		.av_response              (),                                                                      //               (terminated)
		.uav_writeresponserequest (),                                                                      //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                  //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                  //               (terminated)
		.av_writeresponsevalid    ()                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (27),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) flash_ssram_pipeline_bridge_s0_translator (
		.clk                      (pll_c0_out),                                                                                //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                                        //                    reset.reset
		.uav_address              (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (flash_ssram_pipeline_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_chipselect            (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (10),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) slow_peripheral_bridge_s0_translator (
		.clk                      (pll_c0_out),                                                                           //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (slow_peripheral_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_chipselect            (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (27),
		.AV_DATA_W                      (128),
		.UAV_DATA_W                     (128),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (16),
		.UAV_BYTEENABLE_W               (16),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (5),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (16),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_top_clock_bridge_s0_translator (
		.clk                      (pll_c0_out),                                                                          //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (ddr2_top_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) cpu_jtag_debug_module_translator (
		.clk                      (pll_c0_out),                                                                       //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                               //                    reset.reset
		.uav_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (cpu_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (cpu_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (cpu_jtag_debug_module_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (cpu_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (cpu_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (cpu_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (cpu_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_chipselect            (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (27),
		.AV_DATA_W                      (128),
		.UAV_DATA_W                     (128),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (16),
		.UAV_BYTEENABLE_W               (16),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (5),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (16),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_bot_clock_bridge_s0_translator (
		.clk                      (pll_c0_out),                                                                          //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_debugaccess           (ddr2_bot_clock_bridge_s0_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_chipselect            (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dma_0_control_port_slave_translator (
		.clk                      (pll_c0_out),                                                                          //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                                  //                    reset.reset
		.uav_address              (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dma_0_control_port_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dma_0_control_port_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dma_0_control_port_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dma_0_control_port_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dma_0_control_port_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                    //              (terminated)
		.av_begintransfer         (),                                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                                    //              (terminated)
		.av_burstcount            (),                                                                                    //              (terminated)
		.av_byteenable            (),                                                                                    //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                //              (terminated)
		.av_waitrequest           (1'b0),                                                                                //              (terminated)
		.av_writebyteenable       (),                                                                                    //              (terminated)
		.av_lock                  (),                                                                                    //              (terminated)
		.av_clken                 (),                                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                                //              (terminated)
		.av_debugaccess           (),                                                                                    //              (terminated)
		.av_outputenable          (),                                                                                    //              (terminated)
		.uav_response             (),                                                                                    //              (terminated)
		.av_response              (2'b00),                                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                 //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (10),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (10),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) slow_peripheral_bridge_m0_translator (
		.clk                      (pll_c2_out),                                                                   //                       clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                           //                     reset.reset
		.uav_address              (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (slow_peripheral_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (slow_peripheral_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (slow_peripheral_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (slow_peripheral_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read                  (slow_peripheral_bridge_m0_read),                                               //                          .read
		.av_readdata              (slow_peripheral_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (slow_peripheral_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (slow_peripheral_bridge_m0_write),                                              //                          .write
		.av_writedata             (slow_peripheral_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (slow_peripheral_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                         //               (terminated)
		.av_begintransfer         (1'b0),                                                                         //               (terminated)
		.av_chipselect            (1'b0),                                                                         //               (terminated)
		.av_lock                  (1'b0),                                                                         //               (terminated)
		.uav_clken                (),                                                                             //               (terminated)
		.av_clken                 (1'b1),                                                                         //               (terminated)
		.uav_response             (2'b00),                                                                        //               (terminated)
		.av_response              (),                                                                             //               (terminated)
		.uav_writeresponserequest (),                                                                             //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                         //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                         //               (terminated)
		.av_writeresponsevalid    ()                                                                              //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) high_res_timer_s1_translator (
		.clk                      (pll_c2_out),                                                                   //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                           //                    reset.reset
		.uav_address              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (high_res_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (high_res_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (high_res_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (high_res_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (high_res_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                             //              (terminated)
		.av_begintransfer         (),                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                             //              (terminated)
		.av_burstcount            (),                                                                             //              (terminated)
		.av_byteenable            (),                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                             //              (terminated)
		.av_lock                  (),                                                                             //              (terminated)
		.av_clken                 (),                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                         //              (terminated)
		.av_debugaccess           (),                                                                             //              (terminated)
		.av_outputenable          (),                                                                             //              (terminated)
		.uav_response             (),                                                                             //              (terminated)
		.av_response              (2'b00),                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (pll_c2_out),                                                                             //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                     //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) performance_counter_control_slave_translator (
		.clk                      (pll_c2_out),                                                                                   //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                           //                    reset.reset
		.uav_address              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (performance_counter_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (performance_counter_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (performance_counter_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (performance_counter_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (performance_counter_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_read                  (),                                                                                             //              (terminated)
		.av_beginbursttransfer    (),                                                                                             //              (terminated)
		.av_burstcount            (),                                                                                             //              (terminated)
		.av_byteenable            (),                                                                                             //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                         //              (terminated)
		.av_waitrequest           (1'b0),                                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                                             //              (terminated)
		.av_lock                  (),                                                                                             //              (terminated)
		.av_chipselect            (),                                                                                             //              (terminated)
		.av_clken                 (),                                                                                             //              (terminated)
		.uav_clken                (1'b0),                                                                                         //              (terminated)
		.av_debugaccess           (),                                                                                             //              (terminated)
		.av_outputenable          (),                                                                                             //              (terminated)
		.uav_response             (),                                                                                             //              (terminated)
		.av_response              (2'b00),                                                                                        //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                         //              (terminated)
		.uav_writeresponsevalid   (),                                                                                             //              (terminated)
		.av_writeresponserequest  (),                                                                                             //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sys_clk_timer_s1_translator (
		.clk                      (pll_c2_out),                                                                  //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                          //                    reset.reset
		.uav_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sys_clk_timer_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sys_clk_timer_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (sys_clk_timer_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sys_clk_timer_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (sys_clk_timer_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_control_slave_translator (
		.clk                      (pll_c2_out),                                                                     //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                             //                    reset.reset
		.uav_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sysid_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata              (sysid_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write                 (),                                                                               //              (terminated)
		.av_read                  (),                                                                               //              (terminated)
		.av_writedata             (),                                                                               //              (terminated)
		.av_begintransfer         (),                                                                               //              (terminated)
		.av_beginbursttransfer    (),                                                                               //              (terminated)
		.av_burstcount            (),                                                                               //              (terminated)
		.av_byteenable            (),                                                                               //              (terminated)
		.av_readdatavalid         (1'b0),                                                                           //              (terminated)
		.av_waitrequest           (1'b0),                                                                           //              (terminated)
		.av_writebyteenable       (),                                                                               //              (terminated)
		.av_lock                  (),                                                                               //              (terminated)
		.av_chipselect            (),                                                                               //              (terminated)
		.av_clken                 (),                                                                               //              (terminated)
		.uav_clken                (1'b0),                                                                           //              (terminated)
		.av_debugaccess           (),                                                                               //              (terminated)
		.av_outputenable          (),                                                                               //              (terminated)
		.uav_response             (),                                                                               //              (terminated)
		.av_response              (2'b00),                                                                          //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                           //              (terminated)
		.uav_writeresponsevalid   (),                                                                               //              (terminated)
		.av_writeresponserequest  (),                                                                               //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                            //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) fir_dma_control_translator (
		.clk                      (clk),                                                                        //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                         //                    reset.reset
		.uav_address              (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (fir_dma_control_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (fir_dma_control_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (fir_dma_control_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (fir_dma_control_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (fir_dma_control_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (fir_dma_control_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_begintransfer         (),                                                                           //              (terminated)
		.av_beginbursttransfer    (),                                                                           //              (terminated)
		.av_burstcount            (),                                                                           //              (terminated)
		.av_readdatavalid         (1'b0),                                                                       //              (terminated)
		.av_waitrequest           (1'b0),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                           //              (terminated)
		.av_lock                  (),                                                                           //              (terminated)
		.av_chipselect            (),                                                                           //              (terminated)
		.av_clken                 (),                                                                           //              (terminated)
		.uav_clken                (1'b0),                                                                       //              (terminated)
		.av_debugaccess           (),                                                                           //              (terminated)
		.av_outputenable          (),                                                                           //              (terminated)
		.uav_response             (),                                                                           //              (terminated)
		.av_response              (2'b00),                                                                      //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                       //              (terminated)
		.uav_writeresponsevalid   (),                                                                           //              (terminated)
		.av_writeresponserequest  (),                                                                           //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pll_pll_slave_translator (
		.clk                      (clk),                                                                      //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                       //                    reset.reset
		.uav_address              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (pll_pll_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (pll_pll_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (pll_pll_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (pll_pll_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (pll_pll_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_chipselect            (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_pio_s1_translator (
		.clk                      (pll_c2_out),                                                               //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                       //                    reset.reset
		.uav_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (button_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (button_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (button_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (button_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (button_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_pio_s1_translator (
		.clk                      (pll_c2_out),                                                            //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                    //                    reset.reset
		.uav_address              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (15),
		.AV_WRITE_WAIT_CYCLES           (15),
		.AV_SETUP_WAIT_CYCLES           (15),
		.AV_DATA_HOLD_CYCLES            (15)
	) lcd_display_control_slave_translator (
		.clk                      (pll_c2_out),                                                                           //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                   //                    reset.reset
		.uav_address              (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (lcd_display_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (lcd_display_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (lcd_display_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (lcd_display_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (lcd_display_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (lcd_display_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_beginbursttransfer    (),                                                                                     //              (terminated)
		.av_burstcount            (),                                                                                     //              (terminated)
		.av_byteenable            (),                                                                                     //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                 //              (terminated)
		.av_waitrequest           (1'b0),                                                                                 //              (terminated)
		.av_writebyteenable       (),                                                                                     //              (terminated)
		.av_lock                  (),                                                                                     //              (terminated)
		.av_chipselect            (),                                                                                     //              (terminated)
		.av_clken                 (),                                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                                 //              (terminated)
		.av_debugaccess           (),                                                                                     //              (terminated)
		.av_outputenable          (),                                                                                     //              (terminated)
		.uav_response             (),                                                                                     //              (terminated)
		.av_response              (2'b00),                                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (10),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) seven_seg_pio_s1_translator (
		.clk                      (pll_c2_out),                                                                  //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                          //                    reset.reset
		.uav_address              (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (seven_seg_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (seven_seg_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (seven_seg_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (seven_seg_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (seven_seg_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                            //              (terminated)
		.av_begintransfer         (),                                                                            //              (terminated)
		.av_beginbursttransfer    (),                                                                            //              (terminated)
		.av_burstcount            (),                                                                            //              (terminated)
		.av_byteenable            (),                                                                            //              (terminated)
		.av_readdatavalid         (1'b0),                                                                        //              (terminated)
		.av_waitrequest           (1'b0),                                                                        //              (terminated)
		.av_writebyteenable       (),                                                                            //              (terminated)
		.av_lock                  (),                                                                            //              (terminated)
		.av_clken                 (),                                                                            //              (terminated)
		.uav_clken                (1'b0),                                                                        //              (terminated)
		.av_debugaccess           (),                                                                            //              (terminated)
		.av_outputenable          (),                                                                            //              (terminated)
		.uav_response             (),                                                                            //              (terminated)
		.av_response              (2'b00),                                                                       //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                        //              (terminated)
		.uav_writeresponsevalid   (),                                                                            //              (terminated)
		.av_writeresponserequest  (),                                                                            //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                         //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (27),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) flash_ssram_pipeline_bridge_m0_translator (
		.clk                      (pll_c0_out),                                                                        //                       clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                                //                     reset.reset
		.uav_address              (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (flash_ssram_pipeline_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (flash_ssram_pipeline_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (flash_ssram_pipeline_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (flash_ssram_pipeline_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read                  (flash_ssram_pipeline_bridge_m0_read),                                               //                          .read
		.av_readdata              (flash_ssram_pipeline_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (flash_ssram_pipeline_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (flash_ssram_pipeline_bridge_m0_write),                                              //                          .write
		.av_writedata             (flash_ssram_pipeline_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (flash_ssram_pipeline_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                              //               (terminated)
		.av_begintransfer         (1'b0),                                                                              //               (terminated)
		.av_chipselect            (1'b0),                                                                              //               (terminated)
		.av_lock                  (1'b0),                                                                              //               (terminated)
		.uav_clken                (),                                                                                  //               (terminated)
		.av_clken                 (1'b1),                                                                              //               (terminated)
		.uav_response             (2'b00),                                                                             //               (terminated)
		.av_response              (),                                                                                  //               (terminated)
		.uav_writeresponserequest (),                                                                                  //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                              //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                              //               (terminated)
		.av_writeresponsevalid    ()                                                                                   //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (20),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ssram_uas_translator (
		.clk                      (pll_c0_out),                                                           //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                   //                    reset.reset
		.uav_address              (ssram_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ssram_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ssram_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ssram_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ssram_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ssram_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ssram_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (ssram_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ssram_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ssram_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (ssram_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock                  (ssram_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess           (ssram_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                     //              (terminated)
		.av_beginbursttransfer    (),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                     //              (terminated)
		.av_chipselect            (),                                                                     //              (terminated)
		.av_clken                 (),                                                                     //              (terminated)
		.uav_clken                (1'b0),                                                                 //              (terminated)
		.av_outputenable          (),                                                                     //              (terminated)
		.uav_response             (),                                                                     //              (terminated)
		.av_response              (2'b00),                                                                //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                 //              (terminated)
		.uav_writeresponsevalid   (),                                                                     //              (terminated)
		.av_writeresponserequest  (),                                                                     //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                  //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (26),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (2),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (1),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ext_flash_uas_translator (
		.clk                      (pll_c0_out),                                                               //                      clk.clk
		.reset                    (rst_controller_004_reset_out_reset),                                       //                    reset.reset
		.uav_address              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ext_flash_uas_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ext_flash_uas_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ext_flash_uas_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ext_flash_uas_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ext_flash_uas_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount            (ext_flash_uas_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ext_flash_uas_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ext_flash_uas_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (ext_flash_uas_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_lock                  (ext_flash_uas_translator_avalon_anti_slave_0_lock),                        //                         .lock
		.av_debugaccess           (ext_flash_uas_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_chipselect            (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (27),
		.AV_DATA_W                   (128),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (16),
		.UAV_ADDRESS_W               (27),
		.UAV_BURSTCOUNT_W            (5),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (16),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) ddr2_bot_clock_bridge_m0_translator (
		.clk                      (sysclk_bot_out_clk_clk),                                                      //                       clk.clk
		.reset                    (rst_controller_006_reset_out_reset),                                          //                     reset.reset
		.uav_address              (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (ddr2_bot_clock_bridge_m0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (ddr2_bot_clock_bridge_m0_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (ddr2_bot_clock_bridge_m0_burstcount),                                         //                          .burstcount
		.av_byteenable            (ddr2_bot_clock_bridge_m0_byteenable),                                         //                          .byteenable
		.av_read                  (ddr2_bot_clock_bridge_m0_read),                                               //                          .read
		.av_readdata              (ddr2_bot_clock_bridge_m0_readdata),                                           //                          .readdata
		.av_readdatavalid         (ddr2_bot_clock_bridge_m0_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (ddr2_bot_clock_bridge_m0_write),                                              //                          .write
		.av_writedata             (ddr2_bot_clock_bridge_m0_writedata),                                          //                          .writedata
		.av_debugaccess           (ddr2_bot_clock_bridge_m0_debugaccess),                                        //                          .debugaccess
		.av_beginbursttransfer    (1'b0),                                                                        //               (terminated)
		.av_begintransfer         (1'b0),                                                                        //               (terminated)
		.av_chipselect            (1'b0),                                                                        //               (terminated)
		.av_lock                  (1'b0),                                                                        //               (terminated)
		.uav_clken                (),                                                                            //               (terminated)
		.av_clken                 (1'b1),                                                                        //               (terminated)
		.uav_response             (2'b00),                                                                       //               (terminated)
		.av_response              (),                                                                            //               (terminated)
		.uav_writeresponserequest (),                                                                            //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                        //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                        //               (terminated)
		.av_writeresponsevalid    ()                                                                             //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (24),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (3),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (27),
		.UAV_BURSTCOUNT_W               (6),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) ddr2_bot_s1_translator (
		.clk                      (sysclk_bot_out_clk_clk),                                                 //                      clk.clk
		.reset                    (~ddr2_bot_reset_request_n_reset),                                        //                    reset.reset
		.uav_address              (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (ddr2_bot_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (ddr2_bot_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (ddr2_bot_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (ddr2_bot_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (ddr2_bot_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_beginbursttransfer    (ddr2_bot_s1_translator_avalon_anti_slave_0_beginbursttransfer),          //                         .beginbursttransfer
		.av_burstcount            (ddr2_bot_s1_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable            (ddr2_bot_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (ddr2_bot_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (~ddr2_bot_s1_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_begintransfer         (),                                                                       //              (terminated)
		.av_writebyteenable       (),                                                                       //              (terminated)
		.av_lock                  (),                                                                       //              (terminated)
		.av_chipselect            (),                                                                       //              (terminated)
		.av_clken                 (),                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                   //              (terminated)
		.av_debugaccess           (),                                                                       //              (terminated)
		.av_outputenable          (),                                                                       //              (terminated)
		.uav_response             (),                                                                       //              (terminated)
		.av_response              (2'b00),                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                    //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (95),
		.PKT_PROTECTION_L          (93),
		.PKT_BEGIN_BURST           (88),
		.PKT_BURSTWRAP_H           (80),
		.PKT_BURSTWRAP_L           (80),
		.PKT_BURST_SIZE_H          (83),
		.PKT_BURST_SIZE_L          (81),
		.PKT_BURST_TYPE_H          (85),
		.PKT_BURST_TYPE_L          (84),
		.PKT_BYTE_CNT_H            (79),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (90),
		.PKT_SRC_ID_L              (90),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (91),
		.PKT_THREAD_ID_H           (92),
		.PKT_THREAD_ID_L           (92),
		.PKT_CACHE_H               (99),
		.PKT_CACHE_L               (96),
		.PKT_DATA_SIDEBAND_H       (87),
		.PKT_DATA_SIDEBAND_L       (87),
		.PKT_QOS_H                 (89),
		.PKT_QOS_L                 (89),
		.PKT_ADDR_SIDEBAND_H       (86),
		.PKT_ADDR_SIDEBAND_L       (86),
		.PKT_RESPONSE_STATUS_H     (101),
		.PKT_RESPONSE_STATUS_L     (100),
		.ST_DATA_W                 (102),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (5),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fir_dma_write_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk),                                                                              //       clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                               // clk_reset.reset
		.av_address              (fir_dma_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (fir_dma_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (fir_dma_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (fir_dma_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (fir_dma_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (fir_dma_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (fir_dma_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (fir_dma_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (fir_dma_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (fir_dma_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (fir_dma_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (width_adapter_001_src_valid),                                                      //        rp.valid
		.rp_data                 (width_adapter_001_src_data),                                                       //          .data
		.rp_channel              (width_adapter_001_src_channel),                                                    //          .channel
		.rp_startofpacket        (width_adapter_001_src_startofpacket),                                              //          .startofpacket
		.rp_endofpacket          (width_adapter_001_src_endofpacket),                                                //          .endofpacket
		.rp_ready                (width_adapter_001_src_ready),                                                      //          .ready
		.av_response             (),                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (203),
		.PKT_PROTECTION_L          (201),
		.PKT_BEGIN_BURST           (196),
		.PKT_BURSTWRAP_H           (188),
		.PKT_BURSTWRAP_L           (188),
		.PKT_BURST_SIZE_H          (191),
		.PKT_BURST_SIZE_L          (189),
		.PKT_BURST_TYPE_H          (193),
		.PKT_BURST_TYPE_L          (192),
		.PKT_BYTE_CNT_H            (187),
		.PKT_BYTE_CNT_L            (182),
		.PKT_ADDR_H                (175),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (176),
		.PKT_TRANS_POSTED          (177),
		.PKT_TRANS_WRITE           (178),
		.PKT_TRANS_READ            (179),
		.PKT_TRANS_LOCK            (180),
		.PKT_TRANS_EXCLUSIVE       (181),
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_SRC_ID_H              (198),
		.PKT_SRC_ID_L              (198),
		.PKT_DEST_ID_H             (199),
		.PKT_DEST_ID_L             (199),
		.PKT_THREAD_ID_H           (200),
		.PKT_THREAD_ID_L           (200),
		.PKT_CACHE_H               (207),
		.PKT_CACHE_L               (204),
		.PKT_DATA_SIDEBAND_H       (195),
		.PKT_DATA_SIDEBAND_L       (195),
		.PKT_QOS_H                 (197),
		.PKT_QOS_L                 (197),
		.PKT_ADDR_SIDEBAND_H       (194),
		.PKT_ADDR_SIDEBAND_L       (194),
		.PKT_RESPONSE_STATUS_H     (209),
		.PKT_RESPONSE_STATUS_L     (208),
		.ST_DATA_W                 (210),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (5),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk                     (sysclk_top_out_clk_clk),                                                               //       clk.clk
		.reset                   (rst_controller_005_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (width_adapter_003_src_valid),                                                          //        rp.valid
		.rp_data                 (width_adapter_003_src_data),                                                           //          .data
		.rp_channel              (width_adapter_003_src_channel),                                                        //          .channel
		.rp_startofpacket        (width_adapter_003_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket          (width_adapter_003_src_endofpacket),                                                    //          .endofpacket
		.rp_ready                (width_adapter_003_src_ready),                                                          //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (124),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_SRC_ID_H              (126),
		.PKT_SRC_ID_L              (126),
		.PKT_DEST_ID_H             (127),
		.PKT_DEST_ID_L             (127),
		.PKT_BURSTWRAP_H           (116),
		.PKT_BURSTWRAP_L           (116),
		.PKT_BYTE_CNT_H            (115),
		.PKT_BYTE_CNT_L            (110),
		.PKT_PROTECTION_H          (131),
		.PKT_PROTECTION_L          (129),
		.PKT_RESPONSE_STATUS_H     (137),
		.PKT_RESPONSE_STATUS_L     (136),
		.PKT_BURST_SIZE_H          (119),
		.PKT_BURST_SIZE_L          (117),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (138),
		.AVS_BURSTCOUNT_W          (6),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_top_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (sysclk_top_out_clk_clk),                                                           //             clk.clk
		.reset                   (~ddr2_top_reset_request_n_reset),                                                  //       clk_reset.reset
		.m0_address              (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_top_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                           //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                           //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                            //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                   //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                     //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                         //                .channel
		.rf_sink_ready           (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (139),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sysclk_top_out_clk_clk),                                                           //       clk.clk
		.reset             (~ddr2_top_reset_request_n_reset),                                                  // clk_reset.reset
		.in_data           (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (66),
		.FIFO_DEPTH          (128),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (sysclk_top_out_clk_clk),                                                     //       clk.clk
		.reset             (~ddr2_top_reset_request_n_reset),                                            // clk_reset.reset
		.in_data           (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (89),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (79),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.PKT_BURST_TYPE_H          (86),
		.PKT_BURST_TYPE_L          (85),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (88),
		.PKT_DATA_SIDEBAND_L       (88),
		.PKT_QOS_H                 (90),
		.PKT_QOS_L                 (90),
		.PKT_ADDR_SIDEBAND_H       (87),
		.PKT_ADDR_SIDEBAND_L       (87),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (4),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fir_dma_read_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk),                                                                             //       clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                              // clk_reset.reset
		.av_address              (fir_dma_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (fir_dma_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (fir_dma_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (fir_dma_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (fir_dma_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (fir_dma_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (fir_dma_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (fir_dma_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (fir_dma_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (fir_dma_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (fir_dma_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (crosser_003_out_valid),                                                           //        rp.valid
		.rp_data                 (crosser_003_out_data),                                                            //          .data
		.rp_channel              (crosser_003_out_channel),                                                         //          .channel
		.rp_startofpacket        (crosser_003_out_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket          (crosser_003_out_endofpacket),                                                     //          .endofpacket
		.rp_ready                (crosser_003_out_ready),                                                           //          .ready
		.av_response             (),                                                                                // (terminated)
		.av_writeresponserequest (1'b0),                                                                            // (terminated)
		.av_writeresponsevalid   ()                                                                                 // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (89),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (79),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.PKT_BURST_TYPE_H          (86),
		.PKT_BURST_TYPE_L          (85),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (88),
		.PKT_DATA_SIDEBAND_L       (88),
		.PKT_QOS_H                 (90),
		.PKT_QOS_L                 (90),
		.PKT_ADDR_SIDEBAND_H       (87),
		.PKT_ADDR_SIDEBAND_L       (87),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_data_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c0_out),                                                                  //       clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                          // clk_reset.reset
		.av_address              (cpu_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                       //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                        //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                     //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                               //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                 //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                       //          .ready
		.av_response             (),                                                                            // (terminated)
		.av_writeresponserequest (1'b0),                                                                        // (terminated)
		.av_writeresponsevalid   ()                                                                             // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_BEGIN_BURST           (89),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (79),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.PKT_BURST_TYPE_H          (86),
		.PKT_BURST_TYPE_L          (85),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_THREAD_ID_H           (97),
		.PKT_THREAD_ID_L           (97),
		.PKT_CACHE_H               (104),
		.PKT_CACHE_L               (101),
		.PKT_DATA_SIDEBAND_H       (88),
		.PKT_DATA_SIDEBAND_L       (88),
		.PKT_QOS_H                 (90),
		.PKT_QOS_L                 (90),
		.PKT_ADDR_SIDEBAND_H       (87),
		.PKT_ADDR_SIDEBAND_L       (87),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (1),
		.BURSTWRAP_VALUE           (3),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_instruction_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c0_out),                                                                         //       clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                 // clk_reset.reset
		.av_address              (cpu_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (cpu_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (cpu_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (cpu_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (cpu_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (cpu_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (cpu_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (cpu_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (cpu_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (cpu_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_001_rsp_src_valid),                                                          //        rp.valid
		.rp_data                 (limiter_001_rsp_src_data),                                                           //          .data
		.rp_channel              (limiter_001_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket        (limiter_001_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket          (limiter_001_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready                (limiter_001_rsp_src_ready),                                                          //          .ready
		.av_response             (),                                                                                   // (terminated)
		.av_writeresponserequest (1'b0),                                                                               // (terminated)
		.av_writeresponsevalid   ()                                                                                    // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (208),
		.PKT_PROTECTION_L          (206),
		.PKT_BEGIN_BURST           (197),
		.PKT_BURSTWRAP_H           (189),
		.PKT_BURSTWRAP_L           (187),
		.PKT_BURST_SIZE_H          (192),
		.PKT_BURST_SIZE_L          (190),
		.PKT_BURST_TYPE_H          (194),
		.PKT_BURST_TYPE_L          (193),
		.PKT_BYTE_CNT_H            (186),
		.PKT_BYTE_CNT_L            (182),
		.PKT_ADDR_H                (175),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (176),
		.PKT_TRANS_POSTED          (177),
		.PKT_TRANS_WRITE           (178),
		.PKT_TRANS_READ            (179),
		.PKT_TRANS_LOCK            (180),
		.PKT_TRANS_EXCLUSIVE       (181),
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_SRC_ID_H              (201),
		.PKT_SRC_ID_L              (199),
		.PKT_DEST_ID_H             (204),
		.PKT_DEST_ID_L             (202),
		.PKT_THREAD_ID_H           (205),
		.PKT_THREAD_ID_L           (205),
		.PKT_CACHE_H               (212),
		.PKT_CACHE_L               (209),
		.PKT_DATA_SIDEBAND_H       (196),
		.PKT_DATA_SIDEBAND_L       (196),
		.PKT_QOS_H                 (198),
		.PKT_QOS_L                 (198),
		.PKT_ADDR_SIDEBAND_H       (195),
		.PKT_ADDR_SIDEBAND_L       (195),
		.PKT_RESPONSE_STATUS_H     (214),
		.PKT_RESPONSE_STATUS_L     (213),
		.ST_DATA_W                 (215),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (5),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (2),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_read_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c0_out),                                                                    //       clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                            // clk_reset.reset
		.av_address              (dma_0_read_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_0_read_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_0_read_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_0_read_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_0_read_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_0_read_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_0_read_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_0_read_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_0_read_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_0_read_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_0_read_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_003_src2_valid),                                                 //        rp.valid
		.rp_data                 (rsp_xbar_demux_003_src2_data),                                                  //          .data
		.rp_channel              (rsp_xbar_demux_003_src2_channel),                                               //          .channel
		.rp_startofpacket        (rsp_xbar_demux_003_src2_startofpacket),                                         //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_003_src2_endofpacket),                                           //          .endofpacket
		.rp_ready                (rsp_xbar_demux_003_src2_ready),                                                 //          .ready
		.av_response             (),                                                                              // (terminated)
		.av_writeresponserequest (1'b0),                                                                          // (terminated)
		.av_writeresponsevalid   ()                                                                               // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (208),
		.PKT_PROTECTION_L          (206),
		.PKT_BEGIN_BURST           (197),
		.PKT_BURSTWRAP_H           (189),
		.PKT_BURSTWRAP_L           (187),
		.PKT_BURST_SIZE_H          (192),
		.PKT_BURST_SIZE_L          (190),
		.PKT_BURST_TYPE_H          (194),
		.PKT_BURST_TYPE_L          (193),
		.PKT_BYTE_CNT_H            (186),
		.PKT_BYTE_CNT_L            (182),
		.PKT_ADDR_H                (175),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (176),
		.PKT_TRANS_POSTED          (177),
		.PKT_TRANS_WRITE           (178),
		.PKT_TRANS_READ            (179),
		.PKT_TRANS_LOCK            (180),
		.PKT_TRANS_EXCLUSIVE       (181),
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_SRC_ID_H              (201),
		.PKT_SRC_ID_L              (199),
		.PKT_DEST_ID_H             (204),
		.PKT_DEST_ID_L             (202),
		.PKT_THREAD_ID_H           (205),
		.PKT_THREAD_ID_L           (205),
		.PKT_CACHE_H               (212),
		.PKT_CACHE_L               (209),
		.PKT_DATA_SIDEBAND_H       (196),
		.PKT_DATA_SIDEBAND_L       (196),
		.PKT_QOS_H                 (198),
		.PKT_QOS_L                 (198),
		.PKT_ADDR_SIDEBAND_H       (195),
		.PKT_ADDR_SIDEBAND_L       (195),
		.PKT_RESPONSE_STATUS_H     (214),
		.PKT_RESPONSE_STATUS_L     (213),
		.ST_DATA_W                 (215),
		.ST_CHANNEL_W              (6),
		.AV_BURSTCOUNT_W           (5),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (3),
		.BURSTWRAP_VALUE           (7),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_write_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c0_out),                                                                     //       clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                             // clk_reset.reset
		.av_address              (dma_0_write_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (dma_0_write_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (dma_0_write_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (dma_0_write_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (dma_0_write_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (dma_0_write_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (dma_0_write_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (dma_0_write_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (dma_0_write_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (dma_0_write_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (dma_0_write_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_005_src2_valid),                                                  //        rp.valid
		.rp_data                 (rsp_xbar_demux_005_src2_data),                                                   //          .data
		.rp_channel              (rsp_xbar_demux_005_src2_channel),                                                //          .channel
		.rp_startofpacket        (rsp_xbar_demux_005_src2_startofpacket),                                          //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_005_src2_endofpacket),                                            //          .endofpacket
		.rp_ready                (rsp_xbar_demux_005_src2_ready),                                                  //          .ready
		.av_response             (),                                                                               // (terminated)
		.av_writeresponserequest (1'b0),                                                                           // (terminated)
		.av_writeresponsevalid   ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (89),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (79),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                          //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                                  //       clk_reset.reset
		.m0_address              (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                                        //                .channel
		.rf_sink_ready           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                          //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                                  // clk_reset.reset
		.in_data           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                                    //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                                          // (terminated)
		.out_startofpacket (),                                                                                              // (terminated)
		.out_endofpacket   (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (89),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (79),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                     //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src1_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src1_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_003_src1_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src1_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src1_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src1_channel),                                                                //                .channel
		.rf_sink_ready           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (81),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                     //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (128),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                               //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_startofpacket  (1'b0),                                                                                     // (terminated)
		.in_endofpacket    (1'b0),                                                                                     // (terminated)
		.out_startofpacket (),                                                                                         // (terminated)
		.out_endofpacket   (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (197),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_ADDR_H                (175),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (176),
		.PKT_TRANS_POSTED          (177),
		.PKT_TRANS_WRITE           (178),
		.PKT_TRANS_READ            (179),
		.PKT_TRANS_LOCK            (180),
		.PKT_SRC_ID_H              (201),
		.PKT_SRC_ID_L              (199),
		.PKT_DEST_ID_H             (204),
		.PKT_DEST_ID_L             (202),
		.PKT_BURSTWRAP_H           (189),
		.PKT_BURSTWRAP_L           (187),
		.PKT_BYTE_CNT_H            (186),
		.PKT_BYTE_CNT_L            (182),
		.PKT_PROTECTION_H          (208),
		.PKT_PROTECTION_L          (206),
		.PKT_RESPONSE_STATUS_H     (214),
		.PKT_RESPONSE_STATUS_L     (213),
		.PKT_BURST_SIZE_H          (192),
		.PKT_BURST_SIZE_L          (190),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (215),
		.AVS_BURSTCOUNT_W          (5),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                    //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_003_src_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_003_src_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_003_src_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_003_src_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_003_src_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_003_src_channel),                                                                  //                .channel
		.rf_sink_ready           (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (216),
		.FIFO_DEPTH          (73),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                    //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (130),
		.FIFO_DEPTH          (128),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                              //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (89),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (79),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                 //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_004_src_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_mux_004_src_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_mux_004_src_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_mux_004_src_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_004_src_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_mux_004_src_channel),                                                               //                .channel
		.rf_sink_ready           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                 //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                           //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_startofpacket  (1'b0),                                                                                 // (terminated)
		.in_endofpacket    (1'b0),                                                                                 // (terminated)
		.out_startofpacket (),                                                                                     // (terminated)
		.out_endofpacket   (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (197),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_ADDR_H                (175),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (176),
		.PKT_TRANS_POSTED          (177),
		.PKT_TRANS_WRITE           (178),
		.PKT_TRANS_READ            (179),
		.PKT_TRANS_LOCK            (180),
		.PKT_SRC_ID_H              (201),
		.PKT_SRC_ID_L              (199),
		.PKT_DEST_ID_H             (204),
		.PKT_DEST_ID_L             (202),
		.PKT_BURSTWRAP_H           (189),
		.PKT_BURSTWRAP_L           (187),
		.PKT_BYTE_CNT_H            (186),
		.PKT_BYTE_CNT_L            (182),
		.PKT_PROTECTION_H          (208),
		.PKT_PROTECTION_L          (206),
		.PKT_RESPONSE_STATUS_H     (214),
		.PKT_RESPONSE_STATUS_L     (213),
		.PKT_BURST_SIZE_H          (192),
		.PKT_BURST_SIZE_L          (190),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (215),
		.AVS_BURSTCOUNT_W          (5),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                    //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_005_src_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_mux_005_src_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_mux_005_src_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_mux_005_src_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_005_src_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_mux_005_src_channel),                                                                  //                .channel
		.rf_sink_ready           (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (216),
		.FIFO_DEPTH          (73),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                    //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (130),
		.FIFO_DEPTH          (128),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                              //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (89),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (93),
		.PKT_SRC_ID_L              (91),
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_BURSTWRAP_H           (81),
		.PKT_BURSTWRAP_L           (79),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (100),
		.PKT_PROTECTION_L          (98),
		.PKT_RESPONSE_STATUS_H     (106),
		.PKT_RESPONSE_STATUS_L     (105),
		.PKT_BURST_SIZE_H          (84),
		.PKT_BURST_SIZE_L          (82),
		.ST_CHANNEL_W              (6),
		.ST_DATA_W                 (107),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dma_0_control_port_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                                    //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                            //       clk_reset.reset
		.m0_address              (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_003_src5_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_003_src5_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_003_src5_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_003_src5_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_003_src5_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_003_src5_channel),                                                               //                .channel
		.rf_sink_ready           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (108),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                                    //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                            // clk_reset.reset
		.in_data           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                              //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                                    // (terminated)
		.out_startofpacket (),                                                                                        // (terminated)
		.out_endofpacket   (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_BEGIN_BURST           (63),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.PKT_BURST_TYPE_H          (60),
		.PKT_BURST_TYPE_L          (59),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_TRANS_EXCLUSIVE       (51),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_THREAD_ID_H           (73),
		.PKT_THREAD_ID_L           (73),
		.PKT_CACHE_H               (80),
		.PKT_CACHE_L               (77),
		.PKT_DATA_SIDEBAND_H       (62),
		.PKT_DATA_SIDEBAND_L       (62),
		.PKT_QOS_H                 (64),
		.PKT_QOS_L                 (64),
		.PKT_ADDR_SIDEBAND_H       (61),
		.PKT_ADDR_SIDEBAND_L       (61),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (11),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c2_out),                                                                            //       clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.av_address              (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_002_rsp_src_valid),                                                             //        rp.valid
		.rp_data                 (limiter_002_rsp_src_data),                                                              //          .data
		.rp_channel              (limiter_002_rsp_src_channel),                                                           //          .channel
		.rp_startofpacket        (limiter_002_rsp_src_startofpacket),                                                     //          .startofpacket
		.rp_endofpacket          (limiter_002_rsp_src_endofpacket),                                                       //          .endofpacket
		.rp_ready                (limiter_002_rsp_src_ready),                                                             //          .ready
		.av_response             (),                                                                                      // (terminated)
		.av_writeresponserequest (1'b0),                                                                                  // (terminated)
		.av_writeresponsevalid   ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                             //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src0_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src0_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_007_src0_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src0_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src0_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src0_channel),                                                        //                .channel
		.rf_sink_ready           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                             //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                       //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                               //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src1_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src1_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_007_src1_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src1_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src1_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src1_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                       //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                               // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) performance_counter_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                             //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                                     //       clk_reset.reset
		.m0_address              (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src2_ready),                                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src2_valid),                                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_007_src2_data),                                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src2_startofpacket),                                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src2_endofpacket),                                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src2_channel),                                                                        //                .channel
		.rf_sink_ready           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                                  //     (terminated)
		.m0_writeresponserequest (),                                                                                                       //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                    //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                             //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                                     // clk_reset.reset
		.in_data           (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                                   // (terminated)
		.csr_readdata      (),                                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                   // (terminated)
		.almost_full_data  (),                                                                                                       // (terminated)
		.almost_empty_data (),                                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                                   // (terminated)
		.out_empty         (),                                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                                   // (terminated)
		.out_error         (),                                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                                   // (terminated)
		.out_channel       ()                                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                            //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src3_ready),                                                         //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src3_valid),                                                         //                .valid
		.cp_data                 (cmd_xbar_demux_007_src3_data),                                                          //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src3_startofpacket),                                                 //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src3_endofpacket),                                                   //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src3_channel),                                                       //                .channel
		.rf_sink_ready           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                            //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                               //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src4_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src4_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_demux_007_src4_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src4_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src4_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src4_channel),                                                          //                .channel
		.rf_sink_ready           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                    //     (terminated)
		.m0_writeresponserequest (),                                                                                         //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                      //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                               //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                    // (terminated)
		.csr_read          (1'b0),                                                                                     // (terminated)
		.csr_write         (1'b0),                                                                                     // (terminated)
		.csr_readdata      (),                                                                                         // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                     // (terminated)
		.almost_full_data  (),                                                                                         // (terminated)
		.almost_empty_data (),                                                                                         // (terminated)
		.in_empty          (1'b0),                                                                                     // (terminated)
		.out_empty         (),                                                                                         // (terminated)
		.in_error          (1'b0),                                                                                     // (terminated)
		.out_error         (),                                                                                         // (terminated)
		.in_channel        (1'b0),                                                                                     // (terminated)
		.out_channel       ()                                                                                          // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) fir_dma_control_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                  //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (fir_dma_control_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_004_out_ready),                                                                //              cp.ready
		.cp_valid                (crosser_004_out_valid),                                                                //                .valid
		.cp_data                 (crosser_004_out_data),                                                                 //                .data
		.cp_startofpacket        (crosser_004_out_startofpacket),                                                        //                .startofpacket
		.cp_endofpacket          (crosser_004_out_endofpacket),                                                          //                .endofpacket
		.cp_channel              (crosser_004_out_channel),                                                              //                .channel
		.rf_sink_ready           (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                //     (terminated)
		.m0_writeresponserequest (),                                                                                     //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                  //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (fir_dma_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (fir_dma_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk),                                                                            //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                             // clk_reset.reset
		.in_data           (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (fir_dma_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_startofpacket  (1'b0),                                                                           // (terminated)
		.in_endofpacket    (1'b0),                                                                           // (terminated)
		.out_startofpacket (),                                                                               // (terminated)
		.out_endofpacket   (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk),                                                                                //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pll_pll_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (crosser_005_out_ready),                                                              //              cp.ready
		.cp_valid                (crosser_005_out_valid),                                                              //                .valid
		.cp_data                 (crosser_005_out_data),                                                               //                .data
		.cp_startofpacket        (crosser_005_out_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (crosser_005_out_endofpacket),                                                        //                .endofpacket
		.cp_channel              (crosser_005_out_channel),                                                            //                .channel
		.rf_sink_ready           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk),                                                                                //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pll_pll_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk),                                                                          //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                           // clk_reset.reset
		.in_data           (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                         //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src7_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src7_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_007_src7_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src7_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src7_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src7_channel),                                                    //                .channel
		.rf_sink_ready           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                         //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                      //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                              //       clk_reset.reset
		.m0_address              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src8_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src8_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_007_src8_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src8_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src8_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src8_channel),                                                 //                .channel
		.rf_sink_ready           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                      //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                              // clk_reset.reset
		.in_data           (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) lcd_display_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                                     //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                             //       clk_reset.reset
		.m0_address              (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src9_ready),                                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src9_valid),                                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_007_src9_data),                                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src9_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src9_endofpacket),                                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src9_channel),                                                                //                .channel
		.rf_sink_ready           (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                                     //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                          // (terminated)
		.csr_read          (1'b0),                                                                                           // (terminated)
		.csr_write         (1'b0),                                                                                           // (terminated)
		.csr_readdata      (),                                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                           // (terminated)
		.almost_full_data  (),                                                                                               // (terminated)
		.almost_empty_data (),                                                                                               // (terminated)
		.in_empty          (1'b0),                                                                                           // (terminated)
		.out_empty         (),                                                                                               // (terminated)
		.in_error          (1'b0),                                                                                           // (terminated)
		.out_error         (),                                                                                               // (terminated)
		.in_channel        (1'b0),                                                                                           // (terminated)
		.out_channel       ()                                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (63),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (45),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (46),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.PKT_TRANS_READ            (49),
		.PKT_TRANS_LOCK            (50),
		.PKT_SRC_ID_H              (68),
		.PKT_SRC_ID_L              (65),
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_BURSTWRAP_H           (55),
		.PKT_BURSTWRAP_L           (55),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_PROTECTION_H          (76),
		.PKT_PROTECTION_L          (74),
		.PKT_RESPONSE_STATUS_H     (82),
		.PKT_RESPONSE_STATUS_L     (81),
		.PKT_BURST_SIZE_H          (58),
		.PKT_BURST_SIZE_L          (56),
		.ST_CHANNEL_W              (11),
		.ST_DATA_W                 (83),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) seven_seg_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c2_out),                                                                            //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_007_src10_ready),                                                        //              cp.ready
		.cp_valid                (cmd_xbar_demux_007_src10_valid),                                                        //                .valid
		.cp_data                 (cmd_xbar_demux_007_src10_data),                                                         //                .data
		.cp_startofpacket        (cmd_xbar_demux_007_src10_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_007_src10_endofpacket),                                                  //                .endofpacket
		.cp_channel              (cmd_xbar_demux_007_src10_channel),                                                      //                .channel
		.rf_sink_ready           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                 //     (terminated)
		.m0_writeresponserequest (),                                                                                      //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                   //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (84),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c2_out),                                                                            //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_BEGIN_BURST           (80),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.PKT_BURST_TYPE_H          (77),
		.PKT_BURST_TYPE_L          (76),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_TRANS_EXCLUSIVE       (68),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (83),
		.PKT_THREAD_ID_H           (84),
		.PKT_THREAD_ID_L           (84),
		.PKT_CACHE_H               (91),
		.PKT_CACHE_L               (88),
		.PKT_DATA_SIDEBAND_H       (79),
		.PKT_DATA_SIDEBAND_L       (79),
		.PKT_QOS_H                 (81),
		.PKT_QOS_L                 (81),
		.PKT_ADDR_SIDEBAND_H       (78),
		.PKT_ADDR_SIDEBAND_L       (78),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk                     (pll_c0_out),                                                                                 //       clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                         // clk_reset.reset
		.av_address              (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_003_rsp_src_valid),                                                                  //        rp.valid
		.rp_data                 (limiter_003_rsp_src_data),                                                                   //          .data
		.rp_channel              (limiter_003_rsp_src_channel),                                                                //          .channel
		.rp_startofpacket        (limiter_003_rsp_src_startofpacket),                                                          //          .startofpacket
		.rp_endofpacket          (limiter_003_rsp_src_endofpacket),                                                            //          .endofpacket
		.rp_ready                (limiter_003_rsp_src_ready),                                                                  //          .ready
		.av_response             (),                                                                                           // (terminated)
		.av_writeresponserequest (1'b0),                                                                                       // (terminated)
		.av_writeresponsevalid   ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (80),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (62),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (63),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.PKT_TRANS_READ            (66),
		.PKT_TRANS_LOCK            (67),
		.PKT_SRC_ID_H              (82),
		.PKT_SRC_ID_L              (82),
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (83),
		.PKT_BURSTWRAP_H           (72),
		.PKT_BURSTWRAP_L           (72),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_PROTECTION_H          (87),
		.PKT_PROTECTION_L          (85),
		.PKT_RESPONSE_STATUS_H     (93),
		.PKT_RESPONSE_STATUS_L     (92),
		.PKT_BURST_SIZE_H          (75),
		.PKT_BURST_SIZE_L          (73),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (94),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ssram_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                     //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                             //       clk_reset.reset
		.m0_address              (ssram_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ssram_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ssram_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ssram_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ssram_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ssram_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ssram_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ssram_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_008_src0_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_008_src0_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_008_src0_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_008_src0_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_008_src0_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_008_src0_channel),                                                //                .channel
		.rf_sink_ready           (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ssram_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                          //     (terminated)
		.m0_writeresponserequest (),                                                                               //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                            //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (95),
		.FIFO_DEPTH          (6),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                     //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                             // clk_reset.reset
		.in_data           (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ssram_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (62),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_POSTED          (46),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.PKT_TRANS_LOCK            (49),
		.PKT_SRC_ID_H              (64),
		.PKT_SRC_ID_L              (64),
		.PKT_DEST_ID_H             (65),
		.PKT_DEST_ID_L             (65),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (54),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_PROTECTION_H          (69),
		.PKT_PROTECTION_L          (67),
		.PKT_RESPONSE_STATUS_H     (75),
		.PKT_RESPONSE_STATUS_L     (74),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.ST_CHANNEL_W              (2),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_c0_out),                                                                         //             clk.clk
		.reset                   (rst_controller_004_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ext_flash_uas_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                        //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                        //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                         //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                  //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                      //                .channel
		.rf_sink_ready           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_c0_out),                                                                         //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ext_flash_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (4),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_c0_out),                                                                   //       clk.clk
		.reset             (rst_controller_004_reset_out_reset),                                           // clk_reset.reset
		.in_data           (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (198),
		.PKT_PROTECTION_L          (196),
		.PKT_BEGIN_BURST           (191),
		.PKT_BURSTWRAP_H           (183),
		.PKT_BURSTWRAP_L           (183),
		.PKT_BURST_SIZE_H          (186),
		.PKT_BURST_SIZE_L          (184),
		.PKT_BURST_TYPE_H          (188),
		.PKT_BURST_TYPE_L          (187),
		.PKT_BYTE_CNT_H            (182),
		.PKT_BYTE_CNT_L            (177),
		.PKT_ADDR_H                (170),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_COMPRESSED_READ (171),
		.PKT_TRANS_POSTED          (172),
		.PKT_TRANS_WRITE           (173),
		.PKT_TRANS_READ            (174),
		.PKT_TRANS_LOCK            (175),
		.PKT_TRANS_EXCLUSIVE       (176),
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_SRC_ID_H              (193),
		.PKT_SRC_ID_L              (193),
		.PKT_DEST_ID_H             (194),
		.PKT_DEST_ID_L             (194),
		.PKT_THREAD_ID_H           (195),
		.PKT_THREAD_ID_L           (195),
		.PKT_CACHE_H               (202),
		.PKT_CACHE_L               (199),
		.PKT_DATA_SIDEBAND_H       (190),
		.PKT_DATA_SIDEBAND_L       (190),
		.PKT_QOS_H                 (192),
		.PKT_QOS_L                 (192),
		.PKT_ADDR_SIDEBAND_H       (189),
		.PKT_ADDR_SIDEBAND_L       (189),
		.PKT_RESPONSE_STATUS_H     (204),
		.PKT_RESPONSE_STATUS_L     (203),
		.ST_DATA_W                 (205),
		.ST_CHANNEL_W              (1),
		.AV_BURSTCOUNT_W           (5),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent (
		.clk                     (sysclk_bot_out_clk_clk),                                                               //       clk.clk
		.reset                   (rst_controller_006_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (rsp_xbar_demux_020_src0_valid),                                                        //        rp.valid
		.rp_data                 (rsp_xbar_demux_020_src0_data),                                                         //          .data
		.rp_channel              (rsp_xbar_demux_020_src0_channel),                                                      //          .channel
		.rp_startofpacket        (rsp_xbar_demux_020_src0_startofpacket),                                                //          .startofpacket
		.rp_endofpacket          (rsp_xbar_demux_020_src0_endofpacket),                                                  //          .endofpacket
		.rp_ready                (rsp_xbar_demux_020_src0_ready),                                                        //          .ready
		.av_response             (),                                                                                     // (terminated)
		.av_writeresponserequest (1'b0),                                                                                 // (terminated)
		.av_writeresponsevalid   ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (119),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (98),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (99),
		.PKT_TRANS_POSTED          (100),
		.PKT_TRANS_WRITE           (101),
		.PKT_TRANS_READ            (102),
		.PKT_TRANS_LOCK            (103),
		.PKT_SRC_ID_H              (121),
		.PKT_SRC_ID_L              (121),
		.PKT_DEST_ID_H             (122),
		.PKT_DEST_ID_L             (122),
		.PKT_BURSTWRAP_H           (111),
		.PKT_BURSTWRAP_L           (111),
		.PKT_BYTE_CNT_H            (110),
		.PKT_BYTE_CNT_L            (105),
		.PKT_PROTECTION_H          (126),
		.PKT_PROTECTION_L          (124),
		.PKT_RESPONSE_STATUS_H     (132),
		.PKT_RESPONSE_STATUS_L     (131),
		.PKT_BURST_SIZE_H          (114),
		.PKT_BURST_SIZE_L          (112),
		.ST_CHANNEL_W              (1),
		.ST_DATA_W                 (133),
		.AVS_BURSTCOUNT_W          (6),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) ddr2_bot_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (sysclk_bot_out_clk_clk),                                                           //             clk.clk
		.reset                   (~ddr2_bot_reset_request_n_reset),                                                  //       clk_reset.reset
		.m0_address              (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (width_adapter_014_src_ready),                                                      //              cp.ready
		.cp_valid                (width_adapter_014_src_valid),                                                      //                .valid
		.cp_data                 (width_adapter_014_src_data),                                                       //                .data
		.cp_startofpacket        (width_adapter_014_src_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (width_adapter_014_src_endofpacket),                                                //                .endofpacket
		.cp_channel              (width_adapter_014_src_channel),                                                    //                .channel
		.rf_sink_ready           (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (134),
		.FIFO_DEPTH          (33),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (sysclk_bot_out_clk_clk),                                                           //       clk.clk
		.reset             (~ddr2_bot_reset_request_n_reset),                                                  // clk_reset.reset
		.in_data           (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (66),
		.FIFO_DEPTH          (64),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (sysclk_bot_out_clk_clk),                                                     //       clk.clk
		.reset             (~ddr2_bot_reset_request_n_reset),                                            // clk_reset.reset
		.in_data           (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                      // (terminated)
		.csr_read          (1'b0),                                                                       // (terminated)
		.csr_write         (1'b0),                                                                       // (terminated)
		.csr_readdata      (),                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                       // (terminated)
		.almost_full_data  (),                                                                           // (terminated)
		.almost_empty_data (),                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                       // (terminated)
		.out_startofpacket (),                                                                           // (terminated)
		.out_endofpacket   (),                                                                           // (terminated)
		.in_empty          (1'b0),                                                                       // (terminated)
		.out_empty         (),                                                                           // (terminated)
		.in_error          (1'b0),                                                                       // (terminated)
		.out_error         (),                                                                           // (terminated)
		.in_channel        (1'b0),                                                                       // (terminated)
		.out_channel       ()                                                                            // (terminated)
	);

	nios_addr_router addr_router (
		.sink_ready         (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fir_dma_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_src_valid),                                                            //          .valid
		.src_data           (addr_router_src_data),                                                             //          .data
		.src_channel        (addr_router_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                       //          .endofpacket
	);

	nios_addr_router_001 addr_router_001 (
		.sink_ready         (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_top_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sysclk_top_out_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                            //          .valid
		.src_data           (addr_router_001_src_data),                                                             //          .data
		.src_channel        (addr_router_001_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                       //          .endofpacket
	);

	nios_id_router id_router (
		.sink_ready         (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_top_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sysclk_top_out_clk_clk),                                                 //       clk.clk
		.reset              (~ddr2_top_reset_request_n_reset),                                        // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                    //       src.ready
		.src_valid          (id_router_src_valid),                                                    //          .valid
		.src_data           (id_router_src_data),                                                     //          .data
		.src_channel        (id_router_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                               //          .endofpacket
	);

	nios_addr_router_002 addr_router_002 (
		.sink_ready         (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fir_dma_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                             //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                                                       //       src.ready
		.src_valid          (addr_router_002_src_valid),                                                       //          .valid
		.src_data           (addr_router_002_src_data),                                                        //          .data
		.src_channel        (addr_router_002_src_channel),                                                     //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                                                  //          .endofpacket
	);

	nios_addr_router_003 addr_router_003 (
		.sink_ready         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                  //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                                                   //       src.ready
		.src_valid          (addr_router_003_src_valid),                                                   //          .valid
		.src_data           (addr_router_003_src_data),                                                    //          .data
		.src_channel        (addr_router_003_src_channel),                                                 //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                                              //          .endofpacket
	);

	nios_addr_router_004 addr_router_004 (
		.sink_ready         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                         //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_004_src_valid),                                                          //          .valid
		.src_data           (addr_router_004_src_data),                                                           //          .data
		.src_channel        (addr_router_004_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                                                     //          .endofpacket
	);

	nios_addr_router_005 addr_router_005 (
		.sink_ready         (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_read_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                    //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                     //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                     //          .valid
		.src_data           (addr_router_005_src_data),                                                      //          .data
		.src_channel        (addr_router_005_src_channel),                                                   //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                //          .endofpacket
	);

	nios_addr_router_006 addr_router_006 (
		.sink_ready         (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_write_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                     //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (addr_router_006_src_ready),                                                      //       src.ready
		.src_valid          (addr_router_006_src_valid),                                                      //          .valid
		.src_data           (addr_router_006_src_data),                                                       //          .data
		.src_channel        (addr_router_006_src_channel),                                                    //          .channel
		.src_startofpacket  (addr_router_006_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (addr_router_006_src_endofpacket)                                                 //          .endofpacket
	);

	nios_id_router_001 id_router_001 (
		.sink_ready         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (flash_ssram_pipeline_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                                //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                        // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_001_src_valid),                                                                   //          .valid
		.src_data           (id_router_001_src_data),                                                                    //          .data
		.src_channel        (id_router_001_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                              //          .endofpacket
	);

	nios_id_router_002 id_router_002 (
		.sink_ready         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slow_peripheral_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                           //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                              //       src.ready
		.src_valid          (id_router_002_src_valid),                                                              //          .valid
		.src_data           (id_router_002_src_data),                                                               //          .data
		.src_channel        (id_router_002_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                         //          .endofpacket
	);

	nios_id_router_003 id_router_003 (
		.sink_ready         (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_top_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                          //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                                             //          .valid
		.src_data           (id_router_003_src_data),                                                              //          .data
		.src_channel        (id_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	nios_id_router_004 id_router_004 (
		.sink_ready         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (cpu_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                       //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                          //       src.ready
		.src_valid          (id_router_004_src_valid),                                                          //          .valid
		.src_data           (id_router_004_src_data),                                                           //          .data
		.src_channel        (id_router_004_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                                     //          .endofpacket
	);

	nios_id_router_005 id_router_005 (
		.sink_ready         (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_bot_clock_bridge_s0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                          //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                             //       src.ready
		.src_valid          (id_router_005_src_valid),                                                             //          .valid
		.src_data           (id_router_005_src_data),                                                              //          .data
		.src_channel        (id_router_005_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                        //          .endofpacket
	);

	nios_id_router_002 id_router_006 (
		.sink_ready         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dma_0_control_port_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                          //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                             //       src.ready
		.src_valid          (id_router_006_src_valid),                                                             //          .valid
		.src_data           (id_router_006_src_data),                                                              //          .data
		.src_channel        (id_router_006_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                        //          .endofpacket
	);

	nios_addr_router_007 addr_router_007 (
		.sink_ready         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (slow_peripheral_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (addr_router_007_src_ready),                                                             //       src.ready
		.src_valid          (addr_router_007_src_valid),                                                             //          .valid
		.src_data           (addr_router_007_src_data),                                                              //          .data
		.src_channel        (addr_router_007_src_channel),                                                           //          .channel
		.src_startofpacket  (addr_router_007_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (addr_router_007_src_endofpacket)                                                        //          .endofpacket
	);

	nios_id_router_007 id_router_007 (
		.sink_ready         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (high_res_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                   //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                      //       src.ready
		.src_valid          (id_router_007_src_valid),                                                      //          .valid
		.src_data           (id_router_007_src_data),                                                       //          .data
		.src_channel        (id_router_007_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                 //          .endofpacket
	);

	nios_id_router_007 id_router_008 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                             //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                                //       src.ready
		.src_valid          (id_router_008_src_valid),                                                                //          .valid
		.src_data           (id_router_008_src_data),                                                                 //          .data
		.src_channel        (id_router_008_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                           //          .endofpacket
	);

	nios_id_router_007 id_router_009 (
		.sink_ready         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (performance_counter_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                                   //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                           // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                                      //       src.ready
		.src_valid          (id_router_009_src_valid),                                                                      //          .valid
		.src_data           (id_router_009_src_data),                                                                       //          .data
		.src_channel        (id_router_009_src_channel),                                                                    //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                              //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                                 //          .endofpacket
	);

	nios_id_router_007 id_router_010 (
		.sink_ready         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sys_clk_timer_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                                     //       src.ready
		.src_valid          (id_router_010_src_valid),                                                     //          .valid
		.src_data           (id_router_010_src_data),                                                      //          .data
		.src_channel        (id_router_010_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                                //          .endofpacket
	);

	nios_id_router_007 id_router_011 (
		.sink_ready         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                     //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                        //       src.ready
		.src_valid          (id_router_011_src_valid),                                                        //          .valid
		.src_data           (id_router_011_src_data),                                                         //          .data
		.src_channel        (id_router_011_src_channel),                                                      //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                                //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                                   //          .endofpacket
	);

	nios_id_router_007 id_router_012 (
		.sink_ready         (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (fir_dma_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                        //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                    //       src.ready
		.src_valid          (id_router_012_src_valid),                                                    //          .valid
		.src_data           (id_router_012_src_data),                                                     //          .data
		.src_channel        (id_router_012_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                               //          .endofpacket
	);

	nios_id_router_007 id_router_013 (
		.sink_ready         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pll_pll_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk),                                                                      //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                  //       src.ready
		.src_valid          (id_router_013_src_valid),                                                  //          .valid
		.src_data           (id_router_013_src_data),                                                   //          .data
		.src_channel        (id_router_013_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                             //          .endofpacket
	);

	nios_id_router_007 id_router_014 (
		.sink_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                               //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_014_src_ready),                                                  //       src.ready
		.src_valid          (id_router_014_src_valid),                                                  //          .valid
		.src_data           (id_router_014_src_data),                                                   //          .data
		.src_channel        (id_router_014_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_014_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_014_src_endofpacket)                                             //          .endofpacket
	);

	nios_id_router_007 id_router_015 (
		.sink_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                    // clk_reset.reset
		.src_ready          (id_router_015_src_ready),                                               //       src.ready
		.src_valid          (id_router_015_src_valid),                                               //          .valid
		.src_data           (id_router_015_src_data),                                                //          .data
		.src_channel        (id_router_015_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_015_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_015_src_endofpacket)                                          //          .endofpacket
	);

	nios_id_router_007 id_router_016 (
		.sink_ready         (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_display_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (id_router_016_src_ready),                                                              //       src.ready
		.src_valid          (id_router_016_src_valid),                                                              //          .valid
		.src_data           (id_router_016_src_data),                                                               //          .data
		.src_channel        (id_router_016_src_channel),                                                            //          .channel
		.src_startofpacket  (id_router_016_src_startofpacket),                                                      //          .startofpacket
		.src_endofpacket    (id_router_016_src_endofpacket)                                                         //          .endofpacket
	);

	nios_id_router_007 id_router_017 (
		.sink_ready         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (seven_seg_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c2_out),                                                                  //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_017_src_ready),                                                     //       src.ready
		.src_valid          (id_router_017_src_valid),                                                     //          .valid
		.src_data           (id_router_017_src_data),                                                      //          .data
		.src_channel        (id_router_017_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_017_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_017_src_endofpacket)                                                //          .endofpacket
	);

	nios_addr_router_008 addr_router_008 (
		.sink_ready         (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (flash_ssram_pipeline_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                                                 //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (addr_router_008_src_ready),                                                                  //       src.ready
		.src_valid          (addr_router_008_src_valid),                                                                  //          .valid
		.src_data           (addr_router_008_src_data),                                                                   //          .data
		.src_channel        (addr_router_008_src_channel),                                                                //          .channel
		.src_startofpacket  (addr_router_008_src_startofpacket),                                                          //          .startofpacket
		.src_endofpacket    (addr_router_008_src_endofpacket)                                                             //          .endofpacket
	);

	nios_id_router_018 id_router_018 (
		.sink_ready         (ssram_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ssram_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ssram_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ssram_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ssram_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                           //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                   // clk_reset.reset
		.src_ready          (id_router_018_src_ready),                                              //       src.ready
		.src_valid          (id_router_018_src_valid),                                              //          .valid
		.src_data           (id_router_018_src_data),                                               //          .data
		.src_channel        (id_router_018_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_018_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_018_src_endofpacket)                                         //          .endofpacket
	);

	nios_id_router_019 id_router_019 (
		.sink_ready         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ext_flash_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_c0_out),                                                               //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_019_src_ready),                                                  //       src.ready
		.src_valid          (id_router_019_src_valid),                                                  //          .valid
		.src_data           (id_router_019_src_data),                                                   //          .data
		.src_channel        (id_router_019_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_019_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_019_src_endofpacket)                                             //          .endofpacket
	);

	nios_addr_router_009 addr_router_009 (
		.sink_ready         (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_bot_clock_bridge_m0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (sysclk_bot_out_clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_009_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_009_src_valid),                                                            //          .valid
		.src_data           (addr_router_009_src_data),                                                             //          .data
		.src_channel        (addr_router_009_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_009_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_009_src_endofpacket)                                                       //          .endofpacket
	);

	nios_id_router_020 id_router_020 (
		.sink_ready         (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (ddr2_bot_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (sysclk_bot_out_clk_clk),                                                 //       clk.clk
		.reset              (~ddr2_bot_reset_request_n_reset),                                        // clk_reset.reset
		.src_ready          (id_router_020_src_ready),                                                //       src.ready
		.src_valid          (id_router_020_src_valid),                                                //          .valid
		.src_data           (id_router_020_src_data),                                                 //          .data
		.src_channel        (id_router_020_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_020_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_020_src_endofpacket)                                           //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (80),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_004_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_003_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_003_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_003_src_data),           //          .data
		.cmd_sink_channel       (addr_router_003_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_003_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_003_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),              //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),               //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),            //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),      //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),        //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_003_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_003_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_003_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_003_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_003_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_003_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),              //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),              //          .valid
		.rsp_src_data           (limiter_rsp_src_data),               //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),            //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),      //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),        //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)              // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (96),
		.PKT_DEST_ID_L             (94),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (72),
		.PIPELINED                 (0),
		.ST_DATA_W                 (107),
		.ST_CHANNEL_W              (6),
		.VALID_WIDTH               (6),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (78),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_004_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_004_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_004_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_004_src_data),           //          .data
		.cmd_sink_channel       (addr_router_004_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_004_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_004_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_004_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_004_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_004_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_004_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_004_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_004_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (72),
		.PKT_DEST_ID_L             (69),
		.PKT_TRANS_POSTED          (47),
		.PKT_TRANS_WRITE           (48),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (83),
		.ST_CHANNEL_W              (11),
		.VALID_WIDTH               (11),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (54),
		.PKT_BYTE_CNT_L            (52),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (pll_c2_out),                         //       clk.clk
		.reset                  (rst_controller_002_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_007_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_007_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_007_src_data),           //          .data
		.cmd_sink_channel       (addr_router_007_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_007_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_007_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_007_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_007_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_007_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_007_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_007_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_007_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (83),
		.PKT_DEST_ID_L             (83),
		.PKT_TRANS_POSTED          (64),
		.PKT_TRANS_WRITE           (65),
		.MAX_OUTSTANDING_RESPONSES (5),
		.PIPELINED                 (0),
		.ST_DATA_W                 (94),
		.ST_CHANNEL_W              (2),
		.VALID_WIDTH               (2),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (71),
		.PKT_BYTE_CNT_L            (69),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_003 (
		.clk                    (pll_c0_out),                         //       clk.clk
		.reset                  (rst_controller_004_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_008_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_008_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_008_src_data),           //          .data
		.cmd_sink_channel       (addr_router_008_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_008_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_008_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_003_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_003_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_003_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_003_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_003_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_008_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_008_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_008_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_008_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_008_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_008_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_003_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_003_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_003_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_003_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_003_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_003_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_003_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (44),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (62),
		.PKT_BYTE_CNT_H            (53),
		.PKT_BYTE_CNT_L            (51),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (57),
		.PKT_BURST_SIZE_L          (55),
		.PKT_BURST_TYPE_H          (59),
		.PKT_BURST_TYPE_L          (58),
		.PKT_BURSTWRAP_H           (54),
		.PKT_BURSTWRAP_L           (54),
		.PKT_TRANS_COMPRESSED_READ (45),
		.PKT_TRANS_WRITE           (47),
		.PKT_TRANS_READ            (48),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (76),
		.ST_CHANNEL_W              (2),
		.OUT_BYTE_CNT_H            (52),
		.OUT_BURSTWRAP_H           (54),
		.COMPRESSED_READ_SUPPORT   (0),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1),
		.BURSTWRAP_CONST_VALUE     (1)
	) burst_adapter (
		.clk                   (pll_c0_out),                          //       cr0.clk
		.reset                 (rst_controller_004_reset_out_reset),  // cr0_reset.reset
		.sink0_valid           (width_adapter_012_src_valid),         //     sink0.valid
		.sink0_data            (width_adapter_012_src_data),          //          .data
		.sink0_channel         (width_adapter_012_src_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_012_src_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_012_src_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_012_src_ready),         //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (5),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~merged_resets_in_reset_reset_n),   // reset_in0.reset
		.reset_in1  (~merged_resets_in_reset_reset_n),   // reset_in1.reset
		.reset_in2  (~ddr2_top_reset_request_n_reset),   // reset_in2.reset
		.reset_in3  (cpu_jtag_debug_module_reset_reset), // reset_in3.reset
		.reset_in4  (~ddr2_bot_reset_request_n_reset),   // reset_in4.reset
		.clk        (clk_125),                           //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),    // reset_out.reset
		.reset_in5  (1'b0),                              // (terminated)
		.reset_in6  (1'b0),                              // (terminated)
		.reset_in7  (1'b0),                              // (terminated)
		.reset_in8  (1'b0),                              // (terminated)
		.reset_in9  (1'b0),                              // (terminated)
		.reset_in10 (1'b0),                              // (terminated)
		.reset_in11 (1'b0),                              // (terminated)
		.reset_in12 (1'b0),                              // (terminated)
		.reset_in13 (1'b0),                              // (terminated)
		.reset_in14 (1'b0),                              // (terminated)
		.reset_in15 (1'b0)                               // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_001 (
		.reset_in0  (cpu_jtag_debug_module_reset_reset),  // reset_in0.reset
		.clk        (clk_125),                            //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (5),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_002 (
		.reset_in0  (~merged_resets_in_reset_reset_n),    // reset_in0.reset
		.reset_in1  (~merged_resets_in_reset_reset_n),    // reset_in1.reset
		.reset_in2  (~ddr2_top_reset_request_n_reset),    // reset_in2.reset
		.reset_in3  (cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.reset_in4  (~ddr2_bot_reset_request_n_reset),    // reset_in4.reset
		.clk        (pll_c2_out),                         //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (5),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_003 (
		.reset_in0  (~merged_resets_in_reset_reset_n),    // reset_in0.reset
		.reset_in1  (~merged_resets_in_reset_reset_n),    // reset_in1.reset
		.reset_in2  (~ddr2_top_reset_request_n_reset),    // reset_in2.reset
		.reset_in3  (cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.reset_in4  (~ddr2_bot_reset_request_n_reset),    // reset_in4.reset
		.clk        (clk),                                //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (5),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_004 (
		.reset_in0  (~merged_resets_in_reset_reset_n),    // reset_in0.reset
		.reset_in1  (~merged_resets_in_reset_reset_n),    // reset_in1.reset
		.reset_in2  (~ddr2_top_reset_request_n_reset),    // reset_in2.reset
		.reset_in3  (cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.reset_in4  (~ddr2_bot_reset_request_n_reset),    // reset_in4.reset
		.clk        (pll_c0_out),                         //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (5),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_005 (
		.reset_in0  (~merged_resets_in_reset_reset_n),    // reset_in0.reset
		.reset_in1  (~merged_resets_in_reset_reset_n),    // reset_in1.reset
		.reset_in2  (~ddr2_top_reset_request_n_reset),    // reset_in2.reset
		.reset_in3  (cpu_jtag_debug_module_reset_reset),  // reset_in3.reset
		.reset_in4  (~ddr2_bot_reset_request_n_reset),    // reset_in4.reset
		.clk        (sysclk_top_out_clk_clk),             //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (5),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller_006 (
		.reset_in0  (~ddr2_bot_reset_request_n_reset),    // reset_in0.reset
		.reset_in1  (~ddr2_top_reset_request_n_reset),    // reset_in1.reset
		.reset_in2  (~merged_resets_in_reset_reset_n),    // reset_in2.reset
		.reset_in3  (~merged_resets_in_reset_reset_n),    // reset_in3.reset
		.reset_in4  (cpu_jtag_debug_module_reset_reset),  // reset_in4.reset
		.clk        (sysclk_bot_out_clk_clk),             //       clk.clk
		.reset_out  (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	nios_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk),                                //       clk.clk
		.reset              (rst_controller_003_reset_out_reset), // clk_reset.reset
		.sink_ready         (width_adapter_src_ready),            //      sink.ready
		.sink_channel       (width_adapter_src_channel),          //          .channel
		.sink_data          (width_adapter_src_data),             //          .data
		.sink_startofpacket (width_adapter_src_startofpacket),    //          .startofpacket
		.sink_endofpacket   (width_adapter_src_endofpacket),      //          .endofpacket
		.sink_valid         (width_adapter_src_valid),            //          .valid
		.src0_ready         (cmd_xbar_demux_src0_ready),          //      src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),          //          .valid
		.src0_data          (cmd_xbar_demux_src0_data),           //          .data
		.src0_channel       (cmd_xbar_demux_src0_channel),        //          .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket),  //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket)     //          .endofpacket
	);

	nios_cmd_xbar_demux cmd_xbar_demux_001 (
		.clk                (sysclk_top_out_clk_clk),                //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_002_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_002_src_channel),         //          .channel
		.sink_data          (width_adapter_002_src_data),            //          .data
		.sink_startofpacket (width_adapter_002_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_002_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_002_src_valid),           //          .valid
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (sysclk_top_out_clk_clk),                //       clk.clk
		.reset               (~ddr2_top_reset_request_n_reset),       // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (crosser_out_ready),                     //     sink0.ready
		.sink0_valid         (crosser_out_valid),                     //          .valid
		.sink0_channel       (crosser_out_channel),                   //          .channel
		.sink0_data          (crosser_out_data),                      //          .data
		.sink0_startofpacket (crosser_out_startofpacket),             //          .startofpacket
		.sink0_endofpacket   (crosser_out_endofpacket),               //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux rsp_xbar_demux (
		.clk                (sysclk_top_out_clk_clk),            //       clk.clk
		.reset              (~ddr2_top_reset_request_n_reset),   // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_demux_002 cmd_xbar_demux_002 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_002_src_ready),             //      sink.ready
		.sink_channel       (addr_router_002_src_channel),           //          .channel
		.sink_data          (addr_router_002_src_data),              //          .data
		.sink_startofpacket (addr_router_002_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_002_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_002_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_004_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),                 //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),               //           .channel
		.sink_data          (limiter_cmd_src_data),                  //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),         //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),           //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),                // sink_valid.data
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_003_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_003_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_003_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_003_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_003_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_003_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_003_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_003_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_003_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_003_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_003_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_003_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_003_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_003_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_003_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_003_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_003_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_003_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_003_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_003_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_003_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_003_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_003_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_003_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_003_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_003_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_003_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_003_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_003_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_003_src5_endofpacket)    //           .endofpacket
	);

	nios_cmd_xbar_demux_004 cmd_xbar_demux_004 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_004_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_004_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_004_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_004_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_004_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_004_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_004_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_004_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_004_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_004_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_004_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_004_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_004_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_004_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_004_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_004_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_004_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_004_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_004_src3_endofpacket)    //           .endofpacket
	);

	nios_cmd_xbar_demux_005 cmd_xbar_demux_005 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_005_src_ready),             //      sink.ready
		.sink_channel       (addr_router_005_src_channel),           //          .channel
		.sink_data          (addr_router_005_src_data),              //          .data
		.sink_startofpacket (addr_router_005_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_005_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_005_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_demux_005 cmd_xbar_demux_006 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_006_src_ready),             //      sink.ready
		.sink_channel       (addr_router_006_src_channel),           //          .channel
		.sink_data          (addr_router_006_src_data),              //          .data
		.sink_startofpacket (addr_router_006_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_006_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_006_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_mux_001 cmd_xbar_mux_001 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (crosser_002_out_ready),                 //     sink0.ready
		.sink0_valid         (crosser_002_out_valid),                 //          .valid
		.sink0_channel       (crosser_002_out_channel),               //          .channel
		.sink0_data          (crosser_002_out_data),                  //          .data
		.sink0_startofpacket (crosser_002_out_startofpacket),         //          .startofpacket
		.sink0_endofpacket   (crosser_002_out_endofpacket),           //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_004_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_mux_003 cmd_xbar_mux_003 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_004_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_004_src_valid),           //          .valid
		.sink0_channel       (width_adapter_004_src_channel),         //          .channel
		.sink0_data          (width_adapter_004_src_data),            //          .data
		.sink0_startofpacket (width_adapter_004_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_004_src_endofpacket),     //          .endofpacket
		.sink1_ready         (width_adapter_006_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_006_src_valid),           //          .valid
		.sink1_channel       (width_adapter_006_src_channel),         //          .channel
		.sink1_data          (width_adapter_006_src_data),            //          .data
		.sink1_startofpacket (width_adapter_006_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_006_src_endofpacket),     //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_005_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_mux_004 cmd_xbar_mux_004 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src3_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src3_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src3_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src3_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_004_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src2_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_mux_003 cmd_xbar_mux_005 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (width_adapter_005_src_ready),           //     sink0.ready
		.sink0_valid         (width_adapter_005_src_valid),           //          .valid
		.sink0_channel       (width_adapter_005_src_channel),         //          .channel
		.sink0_data          (width_adapter_005_src_data),            //          .data
		.sink0_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink0_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink1_ready         (width_adapter_007_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_007_src_valid),           //          .valid
		.sink1_channel       (width_adapter_007_src_channel),         //          .channel
		.sink1_data          (width_adapter_007_src_data),            //          .data
		.sink1_startofpacket (width_adapter_007_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_007_src_endofpacket),     //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_006_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_006_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_006_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_006_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_001 rsp_xbar_demux_001 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_001_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_001_src2_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_003 rsp_xbar_demux_003 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_003_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_003_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_003_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_003_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_003_src2_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_004 rsp_xbar_demux_004 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_003 rsp_xbar_demux_005 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.src2_ready         (rsp_xbar_demux_005_src2_ready),         //      src2.ready
		.src2_valid         (rsp_xbar_demux_005_src2_valid),         //          .valid
		.src2_data          (rsp_xbar_demux_005_src2_data),          //          .data
		.src2_channel       (rsp_xbar_demux_005_src2_channel),       //          .channel
		.src2_startofpacket (rsp_xbar_demux_005_src2_startofpacket), //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_005_src2_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_mux_003 rsp_xbar_mux_003 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_003_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_003_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (width_adapter_008_src_ready),           //     sink2.ready
		.sink2_valid         (width_adapter_008_src_valid),           //          .valid
		.sink2_channel       (width_adapter_008_src_channel),         //          .channel
		.sink2_data          (width_adapter_008_src_data),            //          .data
		.sink2_startofpacket (width_adapter_008_src_startofpacket),   //          .startofpacket
		.sink2_endofpacket   (width_adapter_008_src_endofpacket),     //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_004_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (width_adapter_010_src_ready),           //     sink4.ready
		.sink4_valid         (width_adapter_010_src_valid),           //          .valid
		.sink4_channel       (width_adapter_010_src_channel),         //          .channel
		.sink4_data          (width_adapter_010_src_data),            //          .data
		.sink4_startofpacket (width_adapter_010_src_startofpacket),   //          .startofpacket
		.sink4_endofpacket   (width_adapter_010_src_endofpacket),     //          .endofpacket
		.sink5_ready         (rsp_xbar_demux_006_src0_ready),         //     sink5.ready
		.sink5_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink5_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink5_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink5_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_mux_004 rsp_xbar_mux_004 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_004_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_004_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_001_src2_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_001_src2_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_001_src2_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_001_src2_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (width_adapter_009_src_ready),           //     sink1.ready
		.sink1_valid         (width_adapter_009_src_valid),           //          .valid
		.sink1_channel       (width_adapter_009_src_channel),         //          .channel
		.sink1_data          (width_adapter_009_src_data),            //          .data
		.sink1_startofpacket (width_adapter_009_src_startofpacket),   //          .startofpacket
		.sink1_endofpacket   (width_adapter_009_src_endofpacket),     //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_004_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (width_adapter_011_src_ready),           //     sink3.ready
		.sink3_valid         (width_adapter_011_src_valid),           //          .valid
		.sink3_channel       (width_adapter_011_src_channel),         //          .channel
		.sink3_data          (width_adapter_011_src_data),            //          .data
		.sink3_startofpacket (width_adapter_011_src_startofpacket),   //          .startofpacket
		.sink3_endofpacket   (width_adapter_011_src_endofpacket)      //          .endofpacket
	);

	nios_cmd_xbar_demux_007 cmd_xbar_demux_007 (
		.clk                 (pll_c2_out),                             //        clk.clk
		.reset               (rst_controller_002_reset_out_reset),     //  clk_reset.reset
		.sink_ready          (limiter_002_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_002_cmd_src_channel),            //           .channel
		.sink_data           (limiter_002_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_002_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_002_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_002_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_007_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_007_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_007_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_007_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_007_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_007_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_007_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_007_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_007_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_007_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_007_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_007_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_007_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_007_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_007_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_007_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_007_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_007_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_007_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_007_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_007_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_007_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_007_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_007_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_007_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_007_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_007_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_007_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_007_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_007_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_007_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_007_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_007_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_007_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_007_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_007_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_007_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_007_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_007_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_007_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_007_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_007_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_007_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_007_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_007_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_007_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_007_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_007_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_007_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_007_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_007_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_007_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_007_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_007_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_007_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_007_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_007_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_007_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_007_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_007_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_007_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_007_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_007_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_007_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_007_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_007_src10_endofpacket)    //           .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_007 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_008 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_009 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_010 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_011 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_012 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_013 (
		.clk                (clk),                                   //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_014 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_014_src_ready),               //      sink.ready
		.sink_channel       (id_router_014_src_channel),             //          .channel
		.sink_data          (id_router_014_src_data),                //          .data
		.sink_startofpacket (id_router_014_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_014_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_014_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_014_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_014_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_014_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_014_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_014_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_015 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_015_src_ready),               //      sink.ready
		.sink_channel       (id_router_015_src_channel),             //          .channel
		.sink_data          (id_router_015_src_data),                //          .data
		.sink_startofpacket (id_router_015_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_015_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_015_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_015_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_015_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_015_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_015_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_015_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_016 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_016_src_ready),               //      sink.ready
		.sink_channel       (id_router_016_src_channel),             //          .channel
		.sink_data          (id_router_016_src_data),                //          .data
		.sink_startofpacket (id_router_016_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_016_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_016_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_016_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_016_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_016_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_016_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_016_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_007 rsp_xbar_demux_017 (
		.clk                (pll_c2_out),                            //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_017_src_ready),               //      sink.ready
		.sink_channel       (id_router_017_src_channel),             //          .channel
		.sink_data          (id_router_017_src_data),                //          .data
		.sink_startofpacket (id_router_017_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_017_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_017_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_017_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_mux_007 rsp_xbar_mux_007 (
		.clk                  (pll_c2_out),                            //       clk.clk
		.reset                (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.src_ready            (rsp_xbar_mux_007_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_007_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_007_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_007_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_007_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_007_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_007_src0_ready),         //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink0_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink0_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink0_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_008_src0_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_009_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_010_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_010_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_011_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_011_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (crosser_006_out_ready),                 //     sink5.ready
		.sink5_valid          (crosser_006_out_valid),                 //          .valid
		.sink5_channel        (crosser_006_out_channel),               //          .channel
		.sink5_data           (crosser_006_out_data),                  //          .data
		.sink5_startofpacket  (crosser_006_out_startofpacket),         //          .startofpacket
		.sink5_endofpacket    (crosser_006_out_endofpacket),           //          .endofpacket
		.sink6_ready          (crosser_007_out_ready),                 //     sink6.ready
		.sink6_valid          (crosser_007_out_valid),                 //          .valid
		.sink6_channel        (crosser_007_out_channel),               //          .channel
		.sink6_data           (crosser_007_out_data),                  //          .data
		.sink6_startofpacket  (crosser_007_out_startofpacket),         //          .startofpacket
		.sink6_endofpacket    (crosser_007_out_endofpacket),           //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_014_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_014_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_014_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_014_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_014_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_014_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_015_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_015_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_015_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_015_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_015_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_015_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_016_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_016_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_016_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_016_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_016_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_016_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_017_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_017_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_017_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_017_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_017_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_017_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_demux_008 cmd_xbar_demux_008 (
		.clk                (pll_c0_out),                            //        clk.clk
		.reset              (rst_controller_004_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_003_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_003_cmd_src_channel),           //           .channel
		.sink_data          (limiter_003_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_003_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_003_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_003_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_008_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_008_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_008_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_008_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_008_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_008_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_008_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_008_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_008_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_008_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_008_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_008_src1_endofpacket)    //           .endofpacket
	);

	nios_rsp_xbar_demux_018 rsp_xbar_demux_018 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_018_src_ready),               //      sink.ready
		.sink_channel       (id_router_018_src_channel),             //          .channel
		.sink_data          (id_router_018_src_data),                //          .data
		.sink_startofpacket (id_router_018_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_018_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_018_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_018_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_demux_018 rsp_xbar_demux_019 (
		.clk                (pll_c0_out),                            //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.sink_ready         (width_adapter_013_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_013_src_channel),         //          .channel
		.sink_data          (width_adapter_013_src_data),            //          .data
		.sink_startofpacket (width_adapter_013_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_013_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_013_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_019_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	nios_rsp_xbar_mux_008 rsp_xbar_mux_008 (
		.clk                 (pll_c0_out),                            //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_008_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_008_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_008_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_008_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_008_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_008_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_018_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_018_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_018_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_018_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_018_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_018_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_019_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_019_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_019_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_019_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_019_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_019_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_demux_009 cmd_xbar_demux_009 (
		.clk                (sysclk_bot_out_clk_clk),                //       clk.clk
		.reset              (rst_controller_006_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_009_src_ready),             //      sink.ready
		.sink_channel       (addr_router_009_src_channel),           //          .channel
		.sink_data          (addr_router_009_src_data),              //          .data
		.sink_startofpacket (addr_router_009_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_009_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_009_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	nios_cmd_xbar_demux_009 rsp_xbar_demux_020 (
		.clk                (sysclk_bot_out_clk_clk),                //       clk.clk
		.reset              (~ddr2_bot_reset_request_n_reset),       // clk_reset.reset
		.sink_ready         (width_adapter_015_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_015_src_channel),         //          .channel
		.sink_data          (width_adapter_015_src_data),            //          .data
		.sink_startofpacket (width_adapter_015_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_015_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_015_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_020_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_020_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_020_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_020_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_020_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_020_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (79),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (80),
		.IN_PKT_BURSTWRAP_L            (80),
		.IN_PKT_BURST_SIZE_H           (83),
		.IN_PKT_BURST_SIZE_L           (81),
		.IN_PKT_RESPONSE_STATUS_H      (101),
		.IN_PKT_RESPONSE_STATUS_L      (100),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (85),
		.IN_PKT_BURST_TYPE_L           (84),
		.IN_ST_DATA_W                  (102),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (115),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (119),
		.OUT_PKT_BURST_SIZE_L          (117),
		.OUT_PKT_RESPONSE_STATUS_H     (137),
		.OUT_PKT_RESPONSE_STATUS_L     (136),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (121),
		.OUT_PKT_BURST_TYPE_L          (120),
		.OUT_ST_DATA_W                 (138),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter (
		.clk                  (clk),                                //       clk.clk
		.reset                (rst_controller_003_reset_out_reset), // clk_reset.reset
		.in_valid             (addr_router_src_valid),              //      sink.valid
		.in_channel           (addr_router_src_channel),            //          .channel
		.in_startofpacket     (addr_router_src_startofpacket),      //          .startofpacket
		.in_endofpacket       (addr_router_src_endofpacket),        //          .endofpacket
		.in_ready             (addr_router_src_ready),              //          .ready
		.in_data              (addr_router_src_data),               //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),      //       src.endofpacket
		.out_data             (width_adapter_src_data),             //          .data
		.out_channel          (width_adapter_src_channel),          //          .channel
		.out_valid            (width_adapter_src_valid),            //          .valid
		.out_ready            (width_adapter_src_ready),            //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),    //          .startofpacket
		.in_command_size_data (3'b000)                              // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (115),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (116),
		.IN_PKT_BURSTWRAP_L            (116),
		.IN_PKT_BURST_SIZE_H           (119),
		.IN_PKT_BURST_SIZE_L           (117),
		.IN_PKT_RESPONSE_STATUS_H      (137),
		.IN_PKT_RESPONSE_STATUS_L      (136),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (121),
		.IN_PKT_BURST_TYPE_L           (120),
		.IN_ST_DATA_W                  (138),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (79),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (83),
		.OUT_PKT_BURST_SIZE_L          (81),
		.OUT_PKT_RESPONSE_STATUS_H     (101),
		.OUT_PKT_RESPONSE_STATUS_L     (100),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (85),
		.OUT_PKT_BURST_TYPE_L          (84),
		.OUT_ST_DATA_W                 (102),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (1)
	) width_adapter_001 (
		.clk                  (clk),                                 //       clk.clk
		.reset                (rst_controller_003_reset_out_reset),  // clk_reset.reset
		.in_valid             (crosser_001_out_valid),               //      sink.valid
		.in_channel           (crosser_001_out_channel),             //          .channel
		.in_startofpacket     (crosser_001_out_startofpacket),       //          .startofpacket
		.in_endofpacket       (crosser_001_out_endofpacket),         //          .endofpacket
		.in_ready             (crosser_001_out_ready),               //          .ready
		.in_data              (crosser_001_out_data),                //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (175),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (187),
		.IN_PKT_BYTE_CNT_L             (182),
		.IN_PKT_TRANS_COMPRESSED_READ  (176),
		.IN_PKT_BURSTWRAP_H            (188),
		.IN_PKT_BURSTWRAP_L            (188),
		.IN_PKT_BURST_SIZE_H           (191),
		.IN_PKT_BURST_SIZE_L           (189),
		.IN_PKT_RESPONSE_STATUS_H      (209),
		.IN_PKT_RESPONSE_STATUS_L      (208),
		.IN_PKT_TRANS_EXCLUSIVE        (181),
		.IN_PKT_BURST_TYPE_H           (193),
		.IN_PKT_BURST_TYPE_L           (192),
		.IN_ST_DATA_W                  (210),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (115),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (119),
		.OUT_PKT_BURST_SIZE_L          (117),
		.OUT_PKT_RESPONSE_STATUS_H     (137),
		.OUT_PKT_RESPONSE_STATUS_L     (136),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (121),
		.OUT_PKT_BURST_TYPE_L          (120),
		.OUT_ST_DATA_W                 (138),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_002 (
		.clk                  (sysclk_top_out_clk_clk),              //       clk.clk
		.reset                (rst_controller_005_reset_out_reset),  // clk_reset.reset
		.in_valid             (addr_router_001_src_valid),           //      sink.valid
		.in_channel           (addr_router_001_src_channel),         //          .channel
		.in_startofpacket     (addr_router_001_src_startofpacket),   //          .startofpacket
		.in_endofpacket       (addr_router_001_src_endofpacket),     //          .endofpacket
		.in_ready             (addr_router_001_src_ready),           //          .ready
		.in_data              (addr_router_001_src_data),            //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (115),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (116),
		.IN_PKT_BURSTWRAP_L            (116),
		.IN_PKT_BURST_SIZE_H           (119),
		.IN_PKT_BURST_SIZE_L           (117),
		.IN_PKT_RESPONSE_STATUS_H      (137),
		.IN_PKT_RESPONSE_STATUS_L      (136),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (121),
		.IN_PKT_BURST_TYPE_L           (120),
		.IN_ST_DATA_W                  (138),
		.OUT_PKT_ADDR_H                (175),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (187),
		.OUT_PKT_BYTE_CNT_L            (182),
		.OUT_PKT_TRANS_COMPRESSED_READ (176),
		.OUT_PKT_BURST_SIZE_H          (191),
		.OUT_PKT_BURST_SIZE_L          (189),
		.OUT_PKT_RESPONSE_STATUS_H     (209),
		.OUT_PKT_RESPONSE_STATUS_L     (208),
		.OUT_PKT_TRANS_EXCLUSIVE       (181),
		.OUT_PKT_BURST_TYPE_H          (193),
		.OUT_PKT_BURST_TYPE_L          (192),
		.OUT_ST_DATA_W                 (210),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_003 (
		.clk                  (sysclk_top_out_clk_clk),              //       clk.clk
		.reset                (rst_controller_005_reset_out_reset),  // clk_reset.reset
		.in_valid             (rsp_xbar_demux_src1_valid),           //      sink.valid
		.in_channel           (rsp_xbar_demux_src1_channel),         //          .channel
		.in_startofpacket     (rsp_xbar_demux_src1_startofpacket),   //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_src1_endofpacket),     //          .endofpacket
		.in_ready             (rsp_xbar_demux_src1_ready),           //          .ready
		.in_data              (rsp_xbar_demux_src1_data),            //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (78),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (81),
		.IN_PKT_BURSTWRAP_L            (79),
		.IN_PKT_BURST_SIZE_H           (84),
		.IN_PKT_BURST_SIZE_L           (82),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (86),
		.IN_PKT_BURST_TYPE_L           (85),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (175),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (186),
		.OUT_PKT_BYTE_CNT_L            (182),
		.OUT_PKT_TRANS_COMPRESSED_READ (176),
		.OUT_PKT_BURST_SIZE_H          (192),
		.OUT_PKT_BURST_SIZE_L          (190),
		.OUT_PKT_RESPONSE_STATUS_H     (214),
		.OUT_PKT_RESPONSE_STATUS_L     (213),
		.OUT_PKT_TRANS_EXCLUSIVE       (181),
		.OUT_PKT_BURST_TYPE_H          (194),
		.OUT_PKT_BURST_TYPE_L          (193),
		.OUT_ST_DATA_W                 (215),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_004 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_003_src2_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_003_src2_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_003_src2_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_003_src2_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_003_src2_ready),         //          .ready
		.in_data              (cmd_xbar_demux_003_src2_data),          //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_004_src_data),            //          .data
		.out_channel          (width_adapter_004_src_channel),         //          .channel
		.out_valid            (width_adapter_004_src_valid),           //          .valid
		.out_ready            (width_adapter_004_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (78),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (81),
		.IN_PKT_BURSTWRAP_L            (79),
		.IN_PKT_BURST_SIZE_H           (84),
		.IN_PKT_BURST_SIZE_L           (82),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (86),
		.IN_PKT_BURST_TYPE_L           (85),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (175),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (186),
		.OUT_PKT_BYTE_CNT_L            (182),
		.OUT_PKT_TRANS_COMPRESSED_READ (176),
		.OUT_PKT_BURST_SIZE_H          (192),
		.OUT_PKT_BURST_SIZE_L          (190),
		.OUT_PKT_RESPONSE_STATUS_H     (214),
		.OUT_PKT_RESPONSE_STATUS_L     (213),
		.OUT_PKT_TRANS_EXCLUSIVE       (181),
		.OUT_PKT_BURST_TYPE_H          (194),
		.OUT_PKT_BURST_TYPE_L          (193),
		.OUT_ST_DATA_W                 (215),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_005 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_003_src4_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_003_src4_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_003_src4_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_003_src4_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_003_src4_ready),         //          .ready
		.in_data              (cmd_xbar_demux_003_src4_data),          //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_005_src_data),            //          .data
		.out_channel          (width_adapter_005_src_channel),         //          .channel
		.out_valid            (width_adapter_005_src_valid),           //          .valid
		.out_ready            (width_adapter_005_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (78),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (81),
		.IN_PKT_BURSTWRAP_L            (79),
		.IN_PKT_BURST_SIZE_H           (84),
		.IN_PKT_BURST_SIZE_L           (82),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (86),
		.IN_PKT_BURST_TYPE_L           (85),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (175),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (186),
		.OUT_PKT_BYTE_CNT_L            (182),
		.OUT_PKT_TRANS_COMPRESSED_READ (176),
		.OUT_PKT_BURST_SIZE_H          (192),
		.OUT_PKT_BURST_SIZE_L          (190),
		.OUT_PKT_RESPONSE_STATUS_H     (214),
		.OUT_PKT_RESPONSE_STATUS_L     (213),
		.OUT_PKT_TRANS_EXCLUSIVE       (181),
		.OUT_PKT_BURST_TYPE_H          (194),
		.OUT_PKT_BURST_TYPE_L          (193),
		.OUT_ST_DATA_W                 (215),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_006 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_004_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_004_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_004_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_004_src1_data),          //          .data
		.out_endofpacket      (width_adapter_006_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_006_src_data),            //          .data
		.out_channel          (width_adapter_006_src_channel),         //          .channel
		.out_valid            (width_adapter_006_src_valid),           //          .valid
		.out_ready            (width_adapter_006_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_006_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (78),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (81),
		.IN_PKT_BURSTWRAP_L            (79),
		.IN_PKT_BURST_SIZE_H           (84),
		.IN_PKT_BURST_SIZE_L           (82),
		.IN_PKT_RESPONSE_STATUS_H      (106),
		.IN_PKT_RESPONSE_STATUS_L      (105),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (86),
		.IN_PKT_BURST_TYPE_L           (85),
		.IN_ST_DATA_W                  (107),
		.OUT_PKT_ADDR_H                (175),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (186),
		.OUT_PKT_BYTE_CNT_L            (182),
		.OUT_PKT_TRANS_COMPRESSED_READ (176),
		.OUT_PKT_BURST_SIZE_H          (192),
		.OUT_PKT_BURST_SIZE_L          (190),
		.OUT_PKT_RESPONSE_STATUS_H     (214),
		.OUT_PKT_RESPONSE_STATUS_L     (213),
		.OUT_PKT_TRANS_EXCLUSIVE       (181),
		.OUT_PKT_BURST_TYPE_H          (194),
		.OUT_PKT_BURST_TYPE_L          (193),
		.OUT_ST_DATA_W                 (215),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_007 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_004_src3_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_004_src3_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_004_src3_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_004_src3_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_004_src3_ready),         //          .ready
		.in_data              (cmd_xbar_demux_004_src3_data),          //          .data
		.out_endofpacket      (width_adapter_007_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_007_src_data),            //          .data
		.out_channel          (width_adapter_007_src_channel),         //          .channel
		.out_valid            (width_adapter_007_src_valid),           //          .valid
		.out_ready            (width_adapter_007_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_007_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (175),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (186),
		.IN_PKT_BYTE_CNT_L             (182),
		.IN_PKT_TRANS_COMPRESSED_READ  (176),
		.IN_PKT_BURSTWRAP_H            (189),
		.IN_PKT_BURSTWRAP_L            (187),
		.IN_PKT_BURST_SIZE_H           (192),
		.IN_PKT_BURST_SIZE_L           (190),
		.IN_PKT_RESPONSE_STATUS_H      (214),
		.IN_PKT_RESPONSE_STATUS_L      (213),
		.IN_PKT_TRANS_EXCLUSIVE        (181),
		.IN_PKT_BURST_TYPE_H           (194),
		.IN_PKT_BURST_TYPE_L           (193),
		.IN_ST_DATA_W                  (215),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (78),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (84),
		.OUT_PKT_BURST_SIZE_L          (82),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (86),
		.OUT_PKT_BURST_TYPE_L          (85),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_008 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_003_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_003_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_003_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_003_src0_data),          //          .data
		.out_endofpacket      (width_adapter_008_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_008_src_data),            //          .data
		.out_channel          (width_adapter_008_src_channel),         //          .channel
		.out_valid            (width_adapter_008_src_valid),           //          .valid
		.out_ready            (width_adapter_008_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_008_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (175),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (186),
		.IN_PKT_BYTE_CNT_L             (182),
		.IN_PKT_TRANS_COMPRESSED_READ  (176),
		.IN_PKT_BURSTWRAP_H            (189),
		.IN_PKT_BURSTWRAP_L            (187),
		.IN_PKT_BURST_SIZE_H           (192),
		.IN_PKT_BURST_SIZE_L           (190),
		.IN_PKT_RESPONSE_STATUS_H      (214),
		.IN_PKT_RESPONSE_STATUS_L      (213),
		.IN_PKT_TRANS_EXCLUSIVE        (181),
		.IN_PKT_BURST_TYPE_H           (194),
		.IN_PKT_BURST_TYPE_L           (193),
		.IN_ST_DATA_W                  (215),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (78),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (84),
		.OUT_PKT_BURST_SIZE_L          (82),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (86),
		.OUT_PKT_BURST_TYPE_L          (85),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_009 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_003_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_003_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_003_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_003_src1_data),          //          .data
		.out_endofpacket      (width_adapter_009_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_009_src_data),            //          .data
		.out_channel          (width_adapter_009_src_channel),         //          .channel
		.out_valid            (width_adapter_009_src_valid),           //          .valid
		.out_ready            (width_adapter_009_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_009_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (175),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (186),
		.IN_PKT_BYTE_CNT_L             (182),
		.IN_PKT_TRANS_COMPRESSED_READ  (176),
		.IN_PKT_BURSTWRAP_H            (189),
		.IN_PKT_BURSTWRAP_L            (187),
		.IN_PKT_BURST_SIZE_H           (192),
		.IN_PKT_BURST_SIZE_L           (190),
		.IN_PKT_RESPONSE_STATUS_H      (214),
		.IN_PKT_RESPONSE_STATUS_L      (213),
		.IN_PKT_TRANS_EXCLUSIVE        (181),
		.IN_PKT_BURST_TYPE_H           (194),
		.IN_PKT_BURST_TYPE_L           (193),
		.IN_ST_DATA_W                  (215),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (78),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (84),
		.OUT_PKT_BURST_SIZE_L          (82),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (86),
		.OUT_PKT_BURST_TYPE_L          (85),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_010 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_005_src0_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_005_src0_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_005_src0_ready),         //          .ready
		.in_data              (rsp_xbar_demux_005_src0_data),          //          .data
		.out_endofpacket      (width_adapter_010_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_010_src_data),            //          .data
		.out_channel          (width_adapter_010_src_channel),         //          .channel
		.out_valid            (width_adapter_010_src_valid),           //          .valid
		.out_ready            (width_adapter_010_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_010_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (175),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (186),
		.IN_PKT_BYTE_CNT_L             (182),
		.IN_PKT_TRANS_COMPRESSED_READ  (176),
		.IN_PKT_BURSTWRAP_H            (189),
		.IN_PKT_BURSTWRAP_L            (187),
		.IN_PKT_BURST_SIZE_H           (192),
		.IN_PKT_BURST_SIZE_L           (190),
		.IN_PKT_RESPONSE_STATUS_H      (214),
		.IN_PKT_RESPONSE_STATUS_L      (213),
		.IN_PKT_TRANS_EXCLUSIVE        (181),
		.IN_PKT_BURST_TYPE_H           (194),
		.IN_PKT_BURST_TYPE_L           (193),
		.IN_ST_DATA_W                  (215),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (78),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (84),
		.OUT_PKT_BURST_SIZE_L          (82),
		.OUT_PKT_RESPONSE_STATUS_H     (106),
		.OUT_PKT_RESPONSE_STATUS_L     (105),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (86),
		.OUT_PKT_BURST_TYPE_L          (85),
		.OUT_ST_DATA_W                 (107),
		.ST_CHANNEL_W                  (6),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_011 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (rsp_xbar_demux_005_src1_valid),         //      sink.valid
		.in_channel           (rsp_xbar_demux_005_src1_channel),       //          .channel
		.in_startofpacket     (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.in_ready             (rsp_xbar_demux_005_src1_ready),         //          .ready
		.in_data              (rsp_xbar_demux_005_src1_data),          //          .data
		.out_endofpacket      (width_adapter_011_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_011_src_data),            //          .data
		.out_channel          (width_adapter_011_src_channel),         //          .channel
		.out_valid            (width_adapter_011_src_valid),           //          .valid
		.out_ready            (width_adapter_011_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_011_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (62),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (71),
		.IN_PKT_BYTE_CNT_L             (69),
		.IN_PKT_TRANS_COMPRESSED_READ  (63),
		.IN_PKT_BURSTWRAP_H            (72),
		.IN_PKT_BURSTWRAP_L            (72),
		.IN_PKT_BURST_SIZE_H           (75),
		.IN_PKT_BURST_SIZE_L           (73),
		.IN_PKT_RESPONSE_STATUS_H      (93),
		.IN_PKT_RESPONSE_STATUS_L      (92),
		.IN_PKT_TRANS_EXCLUSIVE        (68),
		.IN_PKT_BURST_TYPE_H           (77),
		.IN_PKT_BURST_TYPE_L           (76),
		.IN_ST_DATA_W                  (94),
		.OUT_PKT_ADDR_H                (44),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (53),
		.OUT_PKT_BYTE_CNT_L            (51),
		.OUT_PKT_TRANS_COMPRESSED_READ (45),
		.OUT_PKT_BURST_SIZE_H          (57),
		.OUT_PKT_BURST_SIZE_L          (55),
		.OUT_PKT_RESPONSE_STATUS_H     (75),
		.OUT_PKT_RESPONSE_STATUS_L     (74),
		.OUT_PKT_TRANS_EXCLUSIVE       (50),
		.OUT_PKT_BURST_TYPE_H          (59),
		.OUT_PKT_BURST_TYPE_L          (58),
		.OUT_ST_DATA_W                 (76),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_012 (
		.clk                  (pll_c0_out),                            //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_008_src1_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_008_src1_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_008_src1_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_008_src1_ready),         //          .ready
		.in_data              (cmd_xbar_demux_008_src1_data),          //          .data
		.out_endofpacket      (width_adapter_012_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_012_src_data),            //          .data
		.out_channel          (width_adapter_012_src_channel),         //          .channel
		.out_valid            (width_adapter_012_src_valid),           //          .valid
		.out_ready            (width_adapter_012_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_012_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (44),
		.IN_PKT_ADDR_L                 (18),
		.IN_PKT_DATA_H                 (15),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (17),
		.IN_PKT_BYTEEN_L               (16),
		.IN_PKT_BYTE_CNT_H             (53),
		.IN_PKT_BYTE_CNT_L             (51),
		.IN_PKT_TRANS_COMPRESSED_READ  (45),
		.IN_PKT_BURSTWRAP_H            (54),
		.IN_PKT_BURSTWRAP_L            (54),
		.IN_PKT_BURST_SIZE_H           (57),
		.IN_PKT_BURST_SIZE_L           (55),
		.IN_PKT_RESPONSE_STATUS_H      (75),
		.IN_PKT_RESPONSE_STATUS_L      (74),
		.IN_PKT_TRANS_EXCLUSIVE        (50),
		.IN_PKT_BURST_TYPE_H           (59),
		.IN_PKT_BURST_TYPE_L           (58),
		.IN_ST_DATA_W                  (76),
		.OUT_PKT_ADDR_H                (62),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (71),
		.OUT_PKT_BYTE_CNT_L            (69),
		.OUT_PKT_TRANS_COMPRESSED_READ (63),
		.OUT_PKT_BURST_SIZE_H          (75),
		.OUT_PKT_BURST_SIZE_L          (73),
		.OUT_PKT_RESPONSE_STATUS_H     (93),
		.OUT_PKT_RESPONSE_STATUS_L     (92),
		.OUT_PKT_TRANS_EXCLUSIVE       (68),
		.OUT_PKT_BURST_TYPE_H          (77),
		.OUT_PKT_BURST_TYPE_L          (76),
		.OUT_ST_DATA_W                 (94),
		.ST_CHANNEL_W                  (2),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_013 (
		.clk                  (pll_c0_out),                          //       clk.clk
		.reset                (rst_controller_004_reset_out_reset),  // clk_reset.reset
		.in_valid             (id_router_019_src_valid),             //      sink.valid
		.in_channel           (id_router_019_src_channel),           //          .channel
		.in_startofpacket     (id_router_019_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_019_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_019_src_ready),             //          .ready
		.in_data              (id_router_019_src_data),              //          .data
		.out_endofpacket      (width_adapter_013_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_013_src_data),          //          .data
		.out_channel          (width_adapter_013_src_channel),       //          .channel
		.out_valid            (width_adapter_013_src_valid),         //          .valid
		.out_ready            (width_adapter_013_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_013_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (170),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (182),
		.IN_PKT_BYTE_CNT_L             (177),
		.IN_PKT_TRANS_COMPRESSED_READ  (171),
		.IN_PKT_BURSTWRAP_H            (183),
		.IN_PKT_BURSTWRAP_L            (183),
		.IN_PKT_BURST_SIZE_H           (186),
		.IN_PKT_BURST_SIZE_L           (184),
		.IN_PKT_RESPONSE_STATUS_H      (204),
		.IN_PKT_RESPONSE_STATUS_L      (203),
		.IN_PKT_TRANS_EXCLUSIVE        (176),
		.IN_PKT_BURST_TYPE_H           (188),
		.IN_PKT_BURST_TYPE_L           (187),
		.IN_ST_DATA_W                  (205),
		.OUT_PKT_ADDR_H                (98),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (110),
		.OUT_PKT_BYTE_CNT_L            (105),
		.OUT_PKT_TRANS_COMPRESSED_READ (99),
		.OUT_PKT_BURST_SIZE_H          (114),
		.OUT_PKT_BURST_SIZE_L          (112),
		.OUT_PKT_RESPONSE_STATUS_H     (132),
		.OUT_PKT_RESPONSE_STATUS_L     (131),
		.OUT_PKT_TRANS_EXCLUSIVE       (104),
		.OUT_PKT_BURST_TYPE_H          (116),
		.OUT_PKT_BURST_TYPE_L          (115),
		.OUT_ST_DATA_W                 (133),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (0),
		.RESPONSE_PATH                 (0)
	) width_adapter_014 (
		.clk                  (sysclk_bot_out_clk_clk),                //       clk.clk
		.reset                (~ddr2_bot_reset_request_n_reset),       // clk_reset.reset
		.in_valid             (cmd_xbar_demux_009_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_009_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_009_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_009_src0_data),          //          .data
		.out_endofpacket      (width_adapter_014_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_014_src_data),            //          .data
		.out_channel          (width_adapter_014_src_channel),         //          .channel
		.out_valid            (width_adapter_014_src_valid),           //          .valid
		.out_ready            (width_adapter_014_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_014_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                                 // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (98),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (110),
		.IN_PKT_BYTE_CNT_L             (105),
		.IN_PKT_TRANS_COMPRESSED_READ  (99),
		.IN_PKT_BURSTWRAP_H            (111),
		.IN_PKT_BURSTWRAP_L            (111),
		.IN_PKT_BURST_SIZE_H           (114),
		.IN_PKT_BURST_SIZE_L           (112),
		.IN_PKT_RESPONSE_STATUS_H      (132),
		.IN_PKT_RESPONSE_STATUS_L      (131),
		.IN_PKT_TRANS_EXCLUSIVE        (104),
		.IN_PKT_BURST_TYPE_H           (116),
		.IN_PKT_BURST_TYPE_L           (115),
		.IN_ST_DATA_W                  (133),
		.OUT_PKT_ADDR_H                (170),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (182),
		.OUT_PKT_BYTE_CNT_L            (177),
		.OUT_PKT_TRANS_COMPRESSED_READ (171),
		.OUT_PKT_BURST_SIZE_H          (186),
		.OUT_PKT_BURST_SIZE_L          (184),
		.OUT_PKT_RESPONSE_STATUS_H     (204),
		.OUT_PKT_RESPONSE_STATUS_L     (203),
		.OUT_PKT_TRANS_EXCLUSIVE       (176),
		.OUT_PKT_BURST_TYPE_H          (188),
		.OUT_PKT_BURST_TYPE_L          (187),
		.OUT_ST_DATA_W                 (205),
		.ST_CHANNEL_W                  (1),
		.OPTIMIZE_FOR_RSP              (1),
		.RESPONSE_PATH                 (1)
	) width_adapter_015 (
		.clk                  (sysclk_bot_out_clk_clk),              //       clk.clk
		.reset                (~ddr2_bot_reset_request_n_reset),     // clk_reset.reset
		.in_valid             (id_router_020_src_valid),             //      sink.valid
		.in_channel           (id_router_020_src_channel),           //          .channel
		.in_startofpacket     (id_router_020_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_020_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_020_src_ready),             //          .ready
		.in_data              (id_router_020_src_data),              //          .data
		.out_endofpacket      (width_adapter_015_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_015_src_data),          //          .data
		.out_channel          (width_adapter_015_src_channel),       //          .channel
		.out_valid            (width_adapter_015_src_valid),         //          .valid
		.out_ready            (width_adapter_015_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_015_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (138),
		.BITS_PER_SYMBOL     (138),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk),                                //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset), //  in_clk_reset.reset
		.out_clk           (sysclk_top_out_clk_clk),             //       out_clk.clk
		.out_reset         (~ddr2_top_reset_request_n_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (cmd_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (cmd_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (cmd_xbar_demux_src0_channel),        //              .channel
		.in_data           (cmd_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_out_ready),                  //           out.ready
		.out_valid         (crosser_out_valid),                  //              .valid
		.out_startofpacket (crosser_out_startofpacket),          //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),            //              .endofpacket
		.out_channel       (crosser_out_channel),                //              .channel
		.out_data          (crosser_out_data),                   //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (138),
		.BITS_PER_SYMBOL     (138),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (2),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (sysclk_top_out_clk_clk),             //        in_clk.clk
		.in_reset          (~ddr2_top_reset_request_n_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset), // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_src0_ready),          //            in.ready
		.in_valid          (rsp_xbar_demux_src0_valid),          //              .valid
		.in_startofpacket  (rsp_xbar_demux_src0_startofpacket),  //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_src0_endofpacket),    //              .endofpacket
		.in_channel        (rsp_xbar_demux_src0_channel),        //              .channel
		.in_data           (rsp_xbar_demux_src0_data),           //              .data
		.out_ready         (crosser_001_out_ready),              //           out.ready
		.out_valid         (crosser_001_out_valid),              //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),      //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),        //              .endofpacket
		.out_channel       (crosser_001_out_channel),            //              .channel
		.out_data          (crosser_001_out_data),               //              .data
		.in_empty          (1'b0),                               //   (terminated)
		.in_error          (1'b0),                               //   (terminated)
		.out_empty         (),                                   //   (terminated)
		.out_error         ()                                    //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (clk),                                   //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_c0_out),                            //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_002_src0_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_002_src0_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_002_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src0_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_002_src0_channel),       //              .channel
		.in_data           (cmd_xbar_demux_002_src0_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (107),
		.BITS_PER_SYMBOL     (107),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (6),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (pll_c0_out),                            //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                   //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_001_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_001_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_001_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_001_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_001_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_001_src0_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (11),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (pll_c2_out),                            //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                   //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_007_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_007_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_007_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_007_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_007_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_007_src5_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (11),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (pll_c2_out),                            //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk),                                   //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_007_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_007_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_007_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_007_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_007_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_007_src6_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (11),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (clk),                                   //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_c2_out),                            //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_012_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_012_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_012_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_012_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_012_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_012_src0_data),          //              .data
		.out_ready         (crosser_006_out_ready),                 //           out.ready
		.out_valid         (crosser_006_out_valid),                 //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_006_out_channel),               //              .channel
		.out_data          (crosser_006_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (83),
		.BITS_PER_SYMBOL     (83),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (11),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (clk),                                   //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_c2_out),                            //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_013_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_013_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_013_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_013_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_013_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_013_src0_data),          //              .data
		.out_ready         (crosser_007_out_ready),                 //           out.ready
		.out_valid         (crosser_007_out_valid),                 //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_007_out_channel),               //              .channel
		.out_data          (crosser_007_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	nios_irq_mapper irq_mapper (
		.clk           (pll_c0_out),                         //       clk.clk
		.reset         (rst_controller_004_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk),                                //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_004 (
		.receiver_clk   (pll_c2_out),                         //       receiver_clk.clk
		.sender_clk     (pll_c0_out),                         //         sender_clk.clk
		.receiver_reset (rst_controller_002_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_004_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_004_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

endmodule
